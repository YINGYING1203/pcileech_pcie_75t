//
// PCILeech FPGA.
//
// PCIe BAR PIO controller.
//
// The PCILeech BAR PIO controller allows for easy user-implementation on top
// of the PCILeech AXIS128 PCIe TLP streaming interface.
// The controller consists of a read engine and a write engine and pluggable
// user-implemented PCIe BAR implementations (found at bottom of the file).
//
// Considerations:
// - The core handles 1 DWORD read + 1 DWORD write per CLK max. If a lot of
//   data is written / read from the TLP streaming interface the core may
//   drop packet silently.
// - The core reads 1 DWORD of data (without byte enable) per CLK.
// - The core writes 1 DWORD of data (with byte enable) per CLK.
// - All user-implemented cores must have the same latency in CLKs for the
//   returned read data or else undefined behavior will take place.
// - 32-bit addresses are passed for read/writes. Larger BARs than 4GB are
//   not supported due to addressing constraints. Lower bits (LSBs) are the
//   BAR offset, Higher bits (MSBs) are the 32-bit base address of the BAR.
// - DO NOT edit read/write engines.
// - DO edit pcileech_tlps128_bar_controller (to swap bar implementations).
// - DO edit the bar implementations (at bottom of the file, if neccessary).
//
// Example implementations exists below, swap out any of the example cores
// against a core of your use case, or modify existing cores.
// Following test cores exist (see below in this file):
// - pcileech_bar_impl_zerowrite4k = zero-initialized read/write BAR.
//     It's possible to modify contents by use of .coe file.
// - pcileech_bar_impl_loopaddr = test core that loops back the 32-bit
//     address of the current read. Does not support writes.
// - pcileech_bar_impl_none = core without any reply.
// 
// (c) Ulf Frisk, 2024
// Author: Ulf Frisk, pcileech@frizk.net
//

`timescale 1ns / 1ps
`include "pcileech_header.svh"

module pcileech_tlps128_bar_controller(
    input                   rst,
    input                   clk,
    input                   bar_en,
    input [15:0]            pcie_id,
    IfAXIS128.sink_lite     tlps_in,
    IfAXIS128.source        tlps_out
);
    
    // ------------------------------------------------------------------------
    // 1: TLP RECEIVE:
    // Receive incoming BAR requests from the TLP stream:
    // send them onwards to read and write FIFOs
    // ------------------------------------------------------------------------
    wire in_is_wr_ready;
    bit  in_is_wr_last;
    wire in_is_first    = tlps_in.tuser[0];
    wire in_is_bar      = bar_en && (tlps_in.tuser[8:2] != 0);
    wire in_is_rd       = (in_is_first && tlps_in.tlast && ((tlps_in.tdata[31:25] == 7'b0000000) || (tlps_in.tdata[31:25] == 7'b0010000) || (tlps_in.tdata[31:24] == 8'b00000010)));
    wire in_is_wr       = in_is_wr_last || (in_is_first && in_is_wr_ready && ((tlps_in.tdata[31:25] == 7'b0100000) || (tlps_in.tdata[31:25] == 7'b0110000) || (tlps_in.tdata[31:24] == 8'b01000010)));
    
    always @ ( posedge clk )
        if ( rst ) begin
            in_is_wr_last <= 0;
        end
        else if ( tlps_in.tvalid ) begin
            in_is_wr_last <= !tlps_in.tlast && in_is_wr;
        end
    
    wire [6:0]  wr_bar;
    wire [31:0] wr_addr;
    wire [3:0]  wr_be;
    wire [31:0] wr_data;
    wire        wr_valid;
    wire [87:0] rd_req_ctx;
    wire [6:0]  rd_req_bar;
    wire [31:0] rd_req_addr;
    wire        rd_req_valid;
    wire [87:0] rd_rsp_ctx;
    wire [31:0] rd_rsp_data;
    wire        rd_rsp_valid;
        
    pcileech_tlps128_bar_rdengine i_pcileech_tlps128_bar_rdengine(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        // TLPs:
        .pcie_id        ( pcie_id                       ),
        .tlps_in        ( tlps_in                       ),
        .tlps_in_valid  ( tlps_in.tvalid && in_is_bar && in_is_rd ),
        .tlps_out       ( tlps_out                      ),
        // BAR reads:
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_bar     ( rd_req_bar                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid                  ),
        .rd_rsp_ctx     ( rd_rsp_ctx                    ),
        .rd_rsp_data    ( rd_rsp_data                   ),
        .rd_rsp_valid   ( rd_rsp_valid                  )
    );

    pcileech_tlps128_bar_wrengine i_pcileech_tlps128_bar_wrengine(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        // TLPs:
        .tlps_in        ( tlps_in                       ),
        .tlps_in_valid  ( tlps_in.tvalid && in_is_bar && in_is_wr ),
        .tlps_in_ready  ( in_is_wr_ready                ),
        // outgoing BAR writes:
        .wr_bar         ( wr_bar                        ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid                      )
    );
    
    wire [87:0] bar_rsp_ctx[7];
    wire [31:0] bar_rsp_data[7];
    wire        bar_rsp_valid[7];
    
    assign rd_rsp_ctx = bar_rsp_valid[0] ? bar_rsp_ctx[0] :
                        bar_rsp_valid[1] ? bar_rsp_ctx[1] :
                        bar_rsp_valid[2] ? bar_rsp_ctx[2] :
                        bar_rsp_valid[3] ? bar_rsp_ctx[3] :
                        bar_rsp_valid[4] ? bar_rsp_ctx[4] :
                        bar_rsp_valid[5] ? bar_rsp_ctx[5] :
                        bar_rsp_valid[6] ? bar_rsp_ctx[6] : 0;
    assign rd_rsp_data = bar_rsp_valid[0] ? bar_rsp_data[0] :
                        bar_rsp_valid[1] ? bar_rsp_data[1] :
                        bar_rsp_valid[2] ? bar_rsp_data[2] :
                        bar_rsp_valid[3] ? bar_rsp_data[3] :
                        bar_rsp_valid[4] ? bar_rsp_data[4] :
                        bar_rsp_valid[5] ? bar_rsp_data[5] :
                        bar_rsp_valid[6] ? bar_rsp_data[6] : 0;
    assign rd_rsp_valid = bar_rsp_valid[0] || bar_rsp_valid[1] || bar_rsp_valid[2] || bar_rsp_valid[3] || bar_rsp_valid[4] || bar_rsp_valid[5] || bar_rsp_valid[6];
    
     pcileech_bar_impl_bar i_bar0(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[0]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[0] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[0]                ),
        .rd_rsp_data    ( bar_rsp_data[0]               ),
        .rd_rsp_valid   ( bar_rsp_valid[0]              )
    );
    
    pcileech_bar_impl_none i_bar1(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[1]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[1] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[1]                ),
        .rd_rsp_data    ( bar_rsp_data[1]               ),
        .rd_rsp_valid   ( bar_rsp_valid[1]              )
    );
    
    pcileech_bar_impl_none i_bar2(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[2]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[2] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[2]                ),
        .rd_rsp_data    ( bar_rsp_data[2]               ),
        .rd_rsp_valid   ( bar_rsp_valid[2]              )
    );
    
    pcileech_bar_impl_none i_bar3(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[3]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[3] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[3]                ),
        .rd_rsp_data    ( bar_rsp_data[3]               ),
        .rd_rsp_valid   ( bar_rsp_valid[3]              )
    );
    
    pcileech_bar_impl_none i_bar4(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[4]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[4] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[4]                ),
        .rd_rsp_data    ( bar_rsp_data[4]               ),
        .rd_rsp_valid   ( bar_rsp_valid[4]              )
    );
    
    pcileech_bar_impl_none i_bar5(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[5]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[5] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[5]                ),
        .rd_rsp_data    ( bar_rsp_data[5]               ),
        .rd_rsp_valid   ( bar_rsp_valid[5]              )
    );
    
    pcileech_bar_impl_none i_bar6_optrom(
        .rst            ( rst                           ),
        .clk            ( clk                           ),
        .wr_addr        ( wr_addr                       ),
        .wr_be          ( wr_be                         ),
        .wr_data        ( wr_data                       ),
        .wr_valid       ( wr_valid && wr_bar[6]         ),
        .rd_req_ctx     ( rd_req_ctx                    ),
        .rd_req_addr    ( rd_req_addr                   ),
        .rd_req_valid   ( rd_req_valid && rd_req_bar[6] ),
        .rd_rsp_ctx     ( bar_rsp_ctx[6]                ),
        .rd_rsp_data    ( bar_rsp_data[6]               ),
        .rd_rsp_valid   ( bar_rsp_valid[6]              )
    );


endmodule



// ------------------------------------------------------------------------
// BAR WRITE ENGINE:
// Receives BAR WRITE TLPs and output BAR WRITE requests.
// Holds a 2048-byte buffer.
// Input flow rate is 16bytes/CLK (max).
// Output flow rate is 4bytes/CLK.
// If write engine overflows incoming TLP is completely discarded silently.
// ------------------------------------------------------------------------
module pcileech_tlps128_bar_wrengine(
    input                   rst,    
    input                   clk,
    // TLPs:
    IfAXIS128.sink_lite     tlps_in,
    input                   tlps_in_valid,
    output                  tlps_in_ready,
    // outgoing BAR writes:
    output bit [6:0]        wr_bar,
    output bit [31:0]       wr_addr,
    output bit [3:0]        wr_be,
    output bit [31:0]       wr_data,
    output bit              wr_valid
);

    wire            f_rd_en;
    wire [127:0]    f_tdata;
    wire [3:0]      f_tkeepdw;
    wire [8:0]      f_tuser;
    wire            f_tvalid;
    
    bit [127:0]     tdata;
    bit [3:0]       tkeepdw;
    bit             tlast;
    
    bit [3:0]       be_first;
    bit [3:0]       be_last;
    bit             first_dw;
    bit [31:0]      addr;

    fifo_141_141_clk1_bar_wr i_fifo_141_141_clk1_bar_wr(
        .srst           ( rst                           ),
        .clk            ( clk                           ),
        .wr_en          ( tlps_in_valid                 ),
        .din            ( {tlps_in.tuser[8:0], tlps_in.tkeepdw, tlps_in.tdata} ),
        .full           (                               ),
        .prog_empty     ( tlps_in_ready                 ),
        .rd_en          ( f_rd_en                       ),
        .dout           ( {f_tuser, f_tkeepdw, f_tdata} ),    
        .empty          (                               ),
        .valid          ( f_tvalid                      )
    );
    
    // STATE MACHINE:
    `define S_ENGINE_IDLE        3'h0
    `define S_ENGINE_FIRST       3'h1
    `define S_ENGINE_4DW_REQDATA 3'h2
    `define S_ENGINE_TX0         3'h4
    `define S_ENGINE_TX1         3'h5
    `define S_ENGINE_TX2         3'h6
    `define S_ENGINE_TX3         3'h7
    (* KEEP = "TRUE" *) bit [3:0] state = `S_ENGINE_IDLE;
    
    assign f_rd_en = (state == `S_ENGINE_IDLE) ||
                     (state == `S_ENGINE_4DW_REQDATA) ||
                     (state == `S_ENGINE_TX3) ||
                     ((state == `S_ENGINE_TX2 && !tkeepdw[3])) ||
                     ((state == `S_ENGINE_TX1 && !tkeepdw[2])) ||
                     ((state == `S_ENGINE_TX0 && !f_tkeepdw[1]));

    always @ ( posedge clk ) begin
        wr_addr     <= addr;
        wr_valid    <= ((state == `S_ENGINE_TX0) && f_tvalid) || (state == `S_ENGINE_TX1) || (state == `S_ENGINE_TX2) || (state == `S_ENGINE_TX3);
        
    end

    always @ ( posedge clk )
        if ( rst ) begin
            state <= `S_ENGINE_IDLE;
        end
        else case ( state )
            `S_ENGINE_IDLE: begin
                state   <= `S_ENGINE_FIRST;
            end
            `S_ENGINE_FIRST: begin
                if ( f_tvalid && f_tuser[0] ) begin
                    wr_bar      <= f_tuser[8:2];
                    tdata       <= f_tdata;
                    tkeepdw     <= f_tkeepdw;
                    tlast       <= f_tuser[1];
                    first_dw    <= 1;
                    be_first    <= f_tdata[35:32];
                    be_last     <= f_tdata[39:36];
                    if ( f_tdata[31:29] == 8'b010 ) begin       // 3 DW header, with data
                        addr    <= { f_tdata[95:66], 2'b00 };
                        state   <= `S_ENGINE_TX3;
                    end
                    else if ( f_tdata[31:29] == 8'b011 ) begin  // 4 DW header, with data
                        addr    <= { f_tdata[127:98], 2'b00 };
                        state   <= `S_ENGINE_4DW_REQDATA;
                    end 
                end
                else begin
                    state   <= `S_ENGINE_IDLE;
                end
            end 
            `S_ENGINE_4DW_REQDATA: begin
                state   <= `S_ENGINE_TX0;
            end
            `S_ENGINE_TX0: begin
                tdata       <= f_tdata;
                tkeepdw     <= f_tkeepdw;
                tlast       <= f_tuser[1];
                addr        <= addr + 4;
                wr_data     <= { f_tdata[0+00+:8], f_tdata[0+08+:8], f_tdata[0+16+:8], f_tdata[0+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (f_tkeepdw[1] ? 4'hf : be_last);
                state       <= f_tvalid ? (f_tkeepdw[1] ? `S_ENGINE_TX1 : `S_ENGINE_FIRST) : `S_ENGINE_IDLE;
            end
            `S_ENGINE_TX1: begin
                addr        <= addr + 4;
                wr_data     <= { tdata[32+00+:8], tdata[32+08+:8], tdata[32+16+:8], tdata[32+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (tkeepdw[2] ? 4'hf : be_last);
                state       <= tkeepdw[2] ? `S_ENGINE_TX2 : `S_ENGINE_FIRST;
            end
            `S_ENGINE_TX2: begin
                addr        <= addr + 4;
                wr_data     <= { tdata[64+00+:8], tdata[64+08+:8], tdata[64+16+:8], tdata[64+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (tkeepdw[3] ? 4'hf : be_last);
                state       <= tkeepdw[3] ? `S_ENGINE_TX3 : `S_ENGINE_FIRST;
            end
            `S_ENGINE_TX3: begin
                addr        <= addr + 4;
                wr_data     <= { tdata[96+00+:8], tdata[96+08+:8], tdata[96+16+:8], tdata[96+24+:8] };
                first_dw    <= 0;
                wr_be       <= first_dw ? be_first : (!tlast ? 4'hf : be_last);
                state       <= !tlast ? `S_ENGINE_TX0 : `S_ENGINE_FIRST;
            end
        endcase

endmodule



// ------------------------------------------------------------------------
// BAR READ ENGINE:
// Receives BAR READ TLPs and output BAR READ requests.
// ------------------------------------------------------------------------
module pcileech_tlps128_bar_rdengine(
    input                   rst,    
    input                   clk,
    // TLPs:
    input [15:0]            pcie_id,
    IfAXIS128.sink_lite     tlps_in,
    input                   tlps_in_valid,
    IfAXIS128.source        tlps_out,
    // BAR reads:
    output [87:0]           rd_req_ctx,
    output [6:0]            rd_req_bar,
    output [31:0]           rd_req_addr,
    output                  rd_req_valid,
    input  [87:0]           rd_rsp_ctx,
    input  [31:0]           rd_rsp_data,
    input                   rd_rsp_valid
);

    // ------------------------------------------------------------------------
    // 1: PROCESS AND QUEUE INCOMING READ TLPs:
    // ------------------------------------------------------------------------
    wire [10:0] rd1_in_dwlen    = (tlps_in.tdata[9:0] == 0) ? 11'd1024 : {1'b0, tlps_in.tdata[9:0]};
    wire [6:0]  rd1_in_bar      = tlps_in.tuser[8:2];
    wire [15:0] rd1_in_reqid    = tlps_in.tdata[63:48];
    wire [7:0]  rd1_in_tag      = tlps_in.tdata[47:40];
    wire [31:0] rd1_in_addr     = { ((tlps_in.tdata[31:29] == 3'b000) ? tlps_in.tdata[95:66] : tlps_in.tdata[127:98]), 2'b00 };
    wire [73:0] rd1_in_data;
    assign rd1_in_data[73:63]   = rd1_in_dwlen;
    assign rd1_in_data[62:56]   = rd1_in_bar;   
    assign rd1_in_data[55:48]   = rd1_in_tag;
    assign rd1_in_data[47:32]   = rd1_in_reqid;
    assign rd1_in_data[31:0]    = rd1_in_addr;
    
    wire        rd1_out_rden;
    wire [73:0] rd1_out_data;
    wire        rd1_out_valid;
    
    fifo_74_74_clk1_bar_rd1 i_fifo_74_74_clk1_bar_rd1(
        .srst           ( rst                           ),
        .clk            ( clk                           ),
        .wr_en          ( tlps_in_valid                 ),
        .din            ( rd1_in_data                   ),
        .full           (                               ),
        .rd_en          ( rd1_out_rden                  ),
        .dout           ( rd1_out_data                  ),    
        .empty          (                               ),
        .valid          ( rd1_out_valid                 )
    );
    
    // ------------------------------------------------------------------------
    // 2: PROCESS AND SPLIT READ TLPs INTO RESPONSE TLP READ REQUESTS AND QUEUE:
    //    (READ REQUESTS LARGER THAN 128-BYTES WILL BE SPLIT INTO MULTIPLE).
    // ------------------------------------------------------------------------
    
    wire [10:0] rd1_out_dwlen       = rd1_out_data[73:63];
    wire [4:0]  rd1_out_dwlen5      = rd1_out_data[67:63];
    wire [4:0]  rd1_out_addr5       = rd1_out_data[6:2];
    
    // 1st "instant" packet:
    wire [4:0]  rd2_pkt1_dwlen_pre  = ((rd1_out_addr5 + rd1_out_dwlen5 > 6'h20) || ((rd1_out_addr5 != 0) && (rd1_out_dwlen5 == 0))) ? (6'h20 - rd1_out_addr5) : rd1_out_dwlen5;
    wire [5:0]  rd2_pkt1_dwlen      = (rd2_pkt1_dwlen_pre == 0) ? 6'h20 : rd2_pkt1_dwlen_pre;
    wire [10:0] rd2_pkt1_dwlen_next = rd1_out_dwlen - rd2_pkt1_dwlen;
    wire        rd2_pkt1_large      = (rd1_out_dwlen > 32) || (rd1_out_dwlen != rd2_pkt1_dwlen);
    wire        rd2_pkt1_tiny       = (rd1_out_dwlen == 1);
    wire [11:0] rd2_pkt1_bc         = rd1_out_dwlen << 2;
    wire [85:0] rd2_pkt1;
    assign      rd2_pkt1[85:74]     = rd2_pkt1_bc;
    assign      rd2_pkt1[73:63]     = rd2_pkt1_dwlen;
    assign      rd2_pkt1[62:0]      = rd1_out_data[62:0];
    
    // Nth packet (if split should take place):
    bit  [10:0] rd2_total_dwlen;
    wire [10:0] rd2_total_dwlen_next = rd2_total_dwlen - 11'h20;
    
    bit  [85:0] rd2_pkt2;
    wire [10:0] rd2_pkt2_dwlen = rd2_pkt2[73:63];
    wire        rd2_pkt2_large = (rd2_total_dwlen > 11'h20);
    
    wire        rd2_out_rden;
    
    // STATE MACHINE:
    `define S2_ENGINE_REQDATA     1'h0
    `define S2_ENGINE_PROCESSING  1'h1
    (* KEEP = "TRUE" *) bit [0:0] state2 = `S2_ENGINE_REQDATA;
    
    always @ ( posedge clk )
        if ( rst ) begin
            state2 <= `S2_ENGINE_REQDATA;
        end
        else case ( state2 )
            `S2_ENGINE_REQDATA: begin
                if ( rd1_out_valid && rd2_pkt1_large ) begin
                    rd2_total_dwlen <= rd2_pkt1_dwlen_next;                             // dwlen (total remaining)
                    rd2_pkt2[85:74] <= rd2_pkt1_dwlen_next << 2;                        // byte-count
                    rd2_pkt2[73:63] <= (rd2_pkt1_dwlen_next > 11'h20) ? 11'h20 : rd2_pkt1_dwlen_next;   // dwlen next
                    rd2_pkt2[62:12] <= rd1_out_data[62:12];                             // various data
                    rd2_pkt2[11:0]  <= rd1_out_data[11:0] + (rd2_pkt1_dwlen << 2);      // base address (within 4k page)
                    state2 <= `S2_ENGINE_PROCESSING;
                end
            end
            `S2_ENGINE_PROCESSING: begin
                if ( rd2_out_rden ) begin
                    rd2_total_dwlen <= rd2_total_dwlen_next;                                // dwlen (total remaining)
                    rd2_pkt2[85:74] <= rd2_total_dwlen_next << 2;                           // byte-count
                    rd2_pkt2[73:63] <= (rd2_total_dwlen_next > 11'h20) ? 11'h20 : rd2_total_dwlen_next;   // dwlen next
                    rd2_pkt2[62:12] <= rd2_pkt2[62:12];                                     // various data
                    rd2_pkt2[11:0]  <= rd2_pkt2[11:0] + (rd2_pkt2_dwlen << 2);              // base address (within 4k page)
                    if ( !rd2_pkt2_large ) begin
                        state2 <= `S2_ENGINE_REQDATA;
                    end
                end
            end
        endcase
    
    assign rd1_out_rden = rd2_out_rden && (((state2 == `S2_ENGINE_REQDATA) && (!rd1_out_valid || rd2_pkt1_tiny)) || ((state2 == `S2_ENGINE_PROCESSING) && !rd2_pkt2_large));

    wire [85:0] rd2_in_data  = (state2 == `S2_ENGINE_REQDATA) ? rd2_pkt1 : rd2_pkt2;
    wire        rd2_in_valid = rd1_out_valid || ((state2 == `S2_ENGINE_PROCESSING) && rd2_out_rden);

    bit  [85:0] rd2_out_data;
    bit         rd2_out_valid;
    always @ ( posedge clk ) begin
        rd2_out_data    <= rd2_in_valid ? rd2_in_data : rd2_out_data;
        rd2_out_valid   <= rd2_in_valid && !rst;
    end

    // ------------------------------------------------------------------------
    // 3: PROCESS EACH READ REQUEST PACKAGE PER INDIVIDUAL 32-bit READ DWORDS:
    // ------------------------------------------------------------------------

    wire [4:0]  rd2_out_dwlen   = rd2_out_data[67:63];
    wire        rd2_out_last    = (rd2_out_dwlen == 1);
    wire [9:0]  rd2_out_dwaddr  = rd2_out_data[11:2];
    
    wire        rd3_enable;
    
    bit         rd3_process_valid;
    bit         rd3_process_first;
    bit         rd3_process_last;
    bit [4:0]   rd3_process_dwlen;
    bit [9:0]   rd3_process_dwaddr;
    bit [85:0]  rd3_process_data;
    wire        rd3_process_next_last = (rd3_process_dwlen == 2);
    wire        rd3_process_nextnext_last = (rd3_process_dwlen <= 3);
    
    assign rd_req_ctx   = { rd3_process_first, rd3_process_last, rd3_process_data };
    assign rd_req_bar   = rd3_process_data[62:56];
    assign rd_req_addr  = { rd3_process_data[31:12], rd3_process_dwaddr, 2'b00 };
    assign rd_req_valid = rd3_process_valid;
    
    // STATE MACHINE:
    `define S3_ENGINE_REQDATA     1'h0
    `define S3_ENGINE_PROCESSING  1'h1
    (* KEEP = "TRUE" *) bit [0:0] state3 = `S3_ENGINE_REQDATA;
    
    always @ ( posedge clk )
        if ( rst ) begin
            rd3_process_valid   <= 1'b0;
            state3              <= `S3_ENGINE_REQDATA;
        end
        else case ( state3 )
            `S3_ENGINE_REQDATA: begin
                if ( rd2_out_valid ) begin
                    rd3_process_valid       <= 1'b1;
                    rd3_process_first       <= 1'b1;                    // FIRST
                    rd3_process_last        <= rd2_out_last;            // LAST (low 5 bits of dwlen == 1, [max pktlen = 0x20))
                    rd3_process_dwlen       <= rd2_out_dwlen;           // PKT LENGTH IN DW
                    rd3_process_dwaddr      <= rd2_out_dwaddr;          // DWADDR OF THIS DWORD
                    rd3_process_data[85:0]  <= rd2_out_data[85:0];      // FORWARD / SAVE DATA
                    if ( !rd2_out_last ) begin
                        state3 <= `S3_ENGINE_PROCESSING;
                    end
                end
                else begin
                    rd3_process_valid       <= 1'b0;
                end
            end
            `S3_ENGINE_PROCESSING: begin
                rd3_process_first           <= 1'b0;                    // FIRST
                rd3_process_last            <= rd3_process_next_last;   // LAST
                rd3_process_dwlen           <= rd3_process_dwlen - 1;   // LEN DEC
                rd3_process_dwaddr          <= rd3_process_dwaddr + 1;  // ADDR INC
                if ( rd3_process_next_last ) begin
                    state3 <= `S3_ENGINE_REQDATA;
                end
            end
        endcase

    assign rd2_out_rden = rd3_enable && (
        ((state3 == `S3_ENGINE_REQDATA) && (!rd2_out_valid || rd2_out_last)) ||
        ((state3 == `S3_ENGINE_PROCESSING) && rd3_process_nextnext_last));
    
    // ------------------------------------------------------------------------
    // 4: PROCESS RESPONSES:
    // ------------------------------------------------------------------------
    
    wire        rd_rsp_first    = rd_rsp_ctx[87];
    wire        rd_rsp_last     = rd_rsp_ctx[86];
    
    wire [9:0]  rd_rsp_dwlen    = rd_rsp_ctx[72:63];
    wire [11:0] rd_rsp_bc       = rd_rsp_ctx[85:74];
    wire [15:0] rd_rsp_reqid    = rd_rsp_ctx[47:32];
    wire [7:0]  rd_rsp_tag      = rd_rsp_ctx[55:48];
    wire [6:0]  rd_rsp_lowaddr  = rd_rsp_ctx[6:0];
    wire [31:0] rd_rsp_addr     = rd_rsp_ctx[31:0];
    wire [31:0] rd_rsp_data_bs  = { rd_rsp_data[7:0], rd_rsp_data[15:8], rd_rsp_data[23:16], rd_rsp_data[31:24] };
    
    // 1: 32-bit -> 128-bit state machine:
    bit [127:0] tdata;
    bit [3:0]   tkeepdw = 0;
    bit         tlast;
    bit         first   = 1;
    wire        tvalid  = tlast || tkeepdw[3];
    
    always @ ( posedge clk )
        if ( rst ) begin
            tkeepdw <= 0;
            tlast   <= 0;
            first   <= 0;
        end
        else if ( rd_rsp_valid && rd_rsp_first ) begin
            tkeepdw         <= 4'b1111;
            tlast           <= rd_rsp_last;
            first           <= 1'b1;
            tdata[31:0]     <= { 22'b0100101000000000000000, rd_rsp_dwlen };            // format, type, length
            tdata[63:32]    <= { pcie_id[7:0], pcie_id[15:8], 4'b0, rd_rsp_bc };        // pcie_id, byte_count
            tdata[95:64]    <= { rd_rsp_reqid, rd_rsp_tag, 1'b0, rd_rsp_lowaddr };      // req_id, tag, lower_addr
            tdata[127:96]   <= rd_rsp_data_bs;
        end
        else begin
            tlast   <= rd_rsp_valid && rd_rsp_last;
            tkeepdw <= tvalid ? (rd_rsp_valid ? 4'b0001 : 4'b0000) : (rd_rsp_valid ? ((tkeepdw << 1) | 1'b1) : tkeepdw);
            first   <= 0;
            if ( rd_rsp_valid ) begin
                if ( tvalid || !tkeepdw[0] )
                    tdata[31:0]   <= rd_rsp_data_bs;
                if ( !tkeepdw[1] )
                    tdata[63:32]  <= rd_rsp_data_bs;
                if ( !tkeepdw[2] )
                    tdata[95:64]  <= rd_rsp_data_bs;
                if ( !tkeepdw[3] )
                    tdata[127:96] <= rd_rsp_data_bs;   
            end
        end
    
    // 2.1 - submit to output fifo - will feed into mux/pcie core.
    fifo_134_134_clk1_bar_rdrsp i_fifo_134_134_clk1_bar_rdrsp(
        .srst           ( rst                       ),
        .clk            ( clk                       ),
        .din            ( { first, tlast, tkeepdw, tdata } ),
        .wr_en          ( tvalid                    ),
        .rd_en          ( tlps_out.tready           ),
        .dout           ( { tlps_out.tuser[0], tlps_out.tlast, tlps_out.tkeepdw, tlps_out.tdata } ),
        .full           (                           ),
        .empty          (                           ),
        .prog_empty     ( rd3_enable                ),
        .valid          ( tlps_out.tvalid           )
    );
    
    assign tlps_out.tuser[1] = tlps_out.tlast;
    assign tlps_out.tuser[8:2] = 0;
    
    // 2.2 - packet count:
    bit [10:0]  pkt_count       = 0;
    wire        pkt_count_dec   = tlps_out.tvalid && tlps_out.tlast;
    wire        pkt_count_inc   = tvalid && tlast;
    wire [10:0] pkt_count_next  = pkt_count + pkt_count_inc - pkt_count_dec;
    assign tlps_out.has_data    = (pkt_count_next > 0);
    
    always @ ( posedge clk ) begin
        pkt_count <= rst ? 0 : pkt_count_next;
    end

endmodule



// ------------------------------------------------------------------------
// Example BAR implementation that does nothing but drop any read/writes
// silently without generating a response.
// This is only recommended for placeholder designs.
// Latency = N/A.
// ------------------------------------------------------------------------
module pcileech_bar_impl_none(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input  [87:0]       rd_req_ctx,
    input  [31:0]       rd_req_addr,
    input               rd_req_valid,
    // outgoing BAR read replies:
    output bit [87:0]   rd_rsp_ctx,
    output bit [31:0]   rd_rsp_data,
    output bit          rd_rsp_valid
);

    initial rd_rsp_ctx = 0;
    initial rd_rsp_data = 0;
    initial rd_rsp_valid = 0;

endmodule



// ------------------------------------------------------------------------
// Example BAR implementation of "address loopback" which can be useful
// for testing. Any read to a specific BAR address will result in the
// address as response.
// Latency = 2CLKs.
// ------------------------------------------------------------------------
module pcileech_bar_impl_loopaddr(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input [87:0]        rd_req_ctx,
    input [31:0]        rd_req_addr,
    input               rd_req_valid,
    // outgoing BAR read replies:
    output bit [87:0]   rd_rsp_ctx,
    output bit [31:0]   rd_rsp_data,
    output bit          rd_rsp_valid
);

    bit [87:0]      rd_req_ctx_1;
    bit [31:0]      rd_req_addr_1;
    bit             rd_req_valid_1;
    
    always @ ( posedge clk ) begin
        rd_req_ctx_1    <= rd_req_ctx;
        rd_req_addr_1   <= rd_req_addr;
        rd_req_valid_1  <= rd_req_valid;
        rd_rsp_ctx      <= rd_req_ctx_1;
        rd_rsp_data     <= rd_req_addr_1;
        rd_rsp_valid    <= rd_req_valid_1;
    end    

endmodule



// ------------------------------------------------------------------------
// Example BAR implementation of a 4kB writable initial-zero BAR.
// Latency = 2CLKs.
// ------------------------------------------------------------------------
module pcileech_bar_impl_zerowrite4k(
    input               rst,
    input               clk,
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input  [87:0]       rd_req_ctx,
    input  [31:0]       rd_req_addr,
    input               rd_req_valid,
    // outgoing BAR read replies:
    output bit [87:0]   rd_rsp_ctx,
    output bit [31:0]   rd_rsp_data,
    output bit          rd_rsp_valid
);

    bit [87:0]  drd_req_ctx;
    bit         drd_req_valid;
    wire [31:0] doutb;
    
    always @ ( posedge clk ) begin
        drd_req_ctx     <= rd_req_ctx;
        drd_req_valid   <= rd_req_valid;
        rd_rsp_ctx      <= drd_req_ctx;
        rd_rsp_valid    <= drd_req_valid;
        rd_rsp_data     <= doutb; 
    end
    
    bram_bar_zero4k i_bram_bar_zero4k(
        // Port A - write:
        .addra  ( wr_addr[11:2]     ),
        .clka   ( clk               ),
        .dina   ( wr_data           ),
        .ena    ( wr_valid          ),
        .wea    ( wr_be             ),
        // Port A - read (2 CLK latency):
        .addrb  ( rd_req_addr[11:2] ),
        .clkb   ( clk               ),
        .doutb  ( doutb             ),
        .enb    ( rd_req_valid      )
    );

endmodule

/*	{ PROC_THERMAL_MMIO_TJMAX, 0x599c, 16, 0xff },
	{ PROC_THERMAL_MMIO_PP0_TEMP, 0x597c, 0, 0xff },
	{ PROC_THERMAL_MMIO_PP1_TEMP, 0x5980, 0, 0xff },
	{ PROC_THERMAL_MMIO_PKG_TEMP, 0x5978, 0, 0xff },
	{ PROC_THERMAL_MMIO_THRES_0, 0x5820, 8, 0x7F },
	{ PROC_THERMAL_MMIO_THRES_1, 0x5820, 16, 0x7F },
	{ PROC_THERMAL_MMIO_INT_ENABLE_0, 0x5820, 15, 0x01 },
	{ PROC_THERMAL_MMIO_INT_ENABLE_1, 0x5820, 23, 0x01 },
	{ PROC_THERMAL_MMIO_INT_STATUS_0, 0x7200, 6, 0x01 },
	{ PROC_THERMAL_MMIO_INT_STATUS_1, 0x7200, 8, 0x01 },
*/
module pcileech_bar_impl_bar(
    input               rst,
    input               clk,
    // interrupt enable
    // incoming BAR writes:
    input [31:0]        wr_addr,
    input [3:0]         wr_be,
    input [31:0]        wr_data,
    input               wr_valid,
    // incoming BAR reads:
    input  [87:0]       rd_req_ctx,
    input  [31:0]       rd_req_addr,
    input               rd_req_valid,
    // outgoing BAR read replies:
    output reg [87:0]   rd_rsp_ctx,
    output reg [31:0]   rd_rsp_data,
    output reg          rd_rsp_valid
);
                     
    reg [87:0]      drd_req_ctx;
    reg [31:0]      drd_req_addr;
    reg             drd_req_valid;
                  
    reg [31:0]      dwr_addr;
    reg [31:0]      dwr_data;
    reg             dwr_valid;
               
    reg [31:0]      data_32;
    reg [31:0]      tj_max;
    reg [31:0]      pp0_temp;
    reg [31:0]      pp1_temp;
    reg [31:0]      pkg_temp;
    reg [31:0]      thres;
    reg [31:0]      status;
    reg             o_int;
    time number = 0;
    

    always @ (posedge clk) begin
        if (rst) begin
            number <= 0;
            tj_max <= 32'h05640000;
            pp0_temp <= 32'h00000044;
            pkg_temp <= 32'h0000004B;
            pp1_temp <= 32'h00000046;
            status <= 32'h88180242;
        end


        if (((thres >> 15) & 32'h1) &&((status >> 6) & 32'h1) )begin
                o_int <=1;
        end else begin
            o_int <=0;
            status <= 32'h88180242;
            thres <= 32'h809c00;
        end
       

    
        if (pp0_temp != 32'h00000048) begin
            pp0_temp = pp0_temp + 1;
        end else begin
            pp0_temp = 32'h00000044;
        end
        if (pkg_temp != 32'h0000004F) begin
            pkg_temp = pkg_temp + 1;
        end else begin
            pkg_temp = 32'h0000004B;
        end
        if (pp1_temp != 32'h0000004A) begin
            pp1_temp = pp1_temp + 1;
        end else begin
            pp1_temp = 32'h00000046;
        end
        number          <= number + 1;
        drd_req_ctx     <= rd_req_ctx;
        drd_req_valid   <= rd_req_valid;
        dwr_valid       <= wr_valid;
        drd_req_addr    <= rd_req_addr;
        rd_rsp_ctx      <= drd_req_ctx;
        rd_rsp_valid    <= drd_req_valid;
        dwr_addr        <= wr_addr;
        dwr_data        <= wr_data;
        if (drd_req_valid) begin
            case (({drd_req_addr[31:24], drd_req_addr[23:16], drd_req_addr[15:08], drd_req_addr[07:00]}) & 32'hFFFFF)
        32'h599c : rd_rsp_data <= tj_max;
        32'h597c : rd_rsp_data <= pp0_temp;
        32'h5980 : rd_rsp_data <= pp1_temp;
        32'h5978 : rd_rsp_data <= pkg_temp;
        32'h5820 : rd_rsp_data <= thres;
        32'h7200 : rd_rsp_data <= status;
        //16'h0050 : rd_rsp_data <= timer_counter;
        16'h0054 : rd_rsp_data <= o_int;
        //16'h0058 : rd_rsp_data <= status;
        //16'h005c : rd_rsp_data <= thres;
        16'h0060 : rd_rsp_data <= in_rdy;
        16'h0064 : rd_rsp_data <= base_address_register;
        16'h0000 : rd_rsp_data <= 32'h000C0C08;
        16'h0004 : rd_rsp_data <= 32'h0029100C;
        16'h0008 : rd_rsp_data <= 32'h00100C08;
        16'h000C : rd_rsp_data <= 32'h00180C04;
        16'h0010 : rd_rsp_data <= 32'h0021140C;
        16'h0014 : rd_rsp_data <= 32'h001C100C;
        16'h0018 : rd_rsp_data <= 32'h00081410;
        16'h001C : rd_rsp_data <= 32'h00181910;
        16'h0080 : rd_rsp_data <= 32'h10C68000;
        16'h0084 : rd_rsp_data <= 32'hF0F87843;
        16'h0088 : rd_rsp_data <= 32'hFC212480;
        16'h008C : rd_rsp_data <= 32'h0057C001;
        16'h0090 : rd_rsp_data <= 32'h4F9E1000;
        16'h0094 : rd_rsp_data <= 32'h00063C21;
        16'h0098 : rd_rsp_data <= 32'h4FE00000;
        16'h009C : rd_rsp_data <= 32'h0A025B81;
        16'h00A0 : rd_rsp_data <= 32'h9FF0573E;
        16'h00A4 : rd_rsp_data <= 32'h54210FBF;
        16'h00A8 : rd_rsp_data <= 32'h98C011DF;
        16'h00AC : rd_rsp_data <= 32'hA8000000;
        16'h00B0 : rd_rsp_data <= 32'h045E4904;
        16'h00B4 : rd_rsp_data <= 32'h061C003B;
        16'h00B8 : rd_rsp_data <= 32'h8820E21F;
        16'h00BC : rd_rsp_data <= 32'h58155D63;
        16'h00C8 : rd_rsp_data <= 32'h30000000;
        16'h00D4 : rd_rsp_data <= 32'h01041041;
        16'h00D8 : rd_rsp_data <= 32'h08208080;
        16'h00DC : rd_rsp_data <= 32'h1E560820;
        16'h00E0 : rd_rsp_data <= 32'h80627078;
        16'h00E4 : rd_rsp_data <= 32'h504A645D;
        16'h00E8 : rd_rsp_data <= 32'h806C6B68;
        16'h00EC : rd_rsp_data <= 32'h80808080;
        16'h00F0 : rd_rsp_data <= 32'h80808080;
        16'h00F4 : rd_rsp_data <= 32'h0142C3FD;
        16'h00F8 : rd_rsp_data <= 32'h01020FFF;
        16'h00FC : rd_rsp_data <= 32'h01020FFF;
        16'h0100 : rd_rsp_data <= 32'h01020FFF;
        16'h0108 : rd_rsp_data <= 32'h002093C1;
        16'h010C : rd_rsp_data <= 32'h00FFFFFF;
        16'h0110 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0114 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0120 : rd_rsp_data <= 32'h0001D000;
        16'h0128 : rd_rsp_data <= 32'h03800000;
        16'h012C : rd_rsp_data <= 32'h07458BBC;
        16'h013C : rd_rsp_data <= 32'h023404E3;
        16'h0140 : rd_rsp_data <= 32'h0006087E;
        16'h0148 : rd_rsp_data <= 32'h80100010;
        16'h014C : rd_rsp_data <= 32'h99999999;
        16'h0150 : rd_rsp_data <= 32'h21084210;
        16'h0154 : rd_rsp_data <= 32'h21084210;
        16'h0158 : rd_rsp_data <= 32'h210841F0;
        16'h015C : rd_rsp_data <= 32'h21084210;
        16'h0160 : rd_rsp_data <= 32'h21084270;
        16'h0164 : rd_rsp_data <= 32'h21084270;
        16'h0168 : rd_rsp_data <= 32'h21084250;
        16'h016C : rd_rsp_data <= 32'h21084270;
        16'h0170 : rd_rsp_data <= 32'h21084210;
        16'h0174 : rd_rsp_data <= 32'h21084210;
        16'h0178 : rd_rsp_data <= 32'h00084210;
        16'h017C : rd_rsp_data <= 32'h00077054;
        16'h0180 : rd_rsp_data <= 32'h08400000;
        16'h0198 : rd_rsp_data <= 32'h808CF60A;
        16'h019C : rd_rsp_data <= 32'h00000016;
        16'h01A0 : rd_rsp_data <= 32'h00019400;
        16'h01AC : rd_rsp_data <= 32'h03260244;
        16'h01B0 : rd_rsp_data <= 32'h12481000;
        16'h01B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h01B8 : rd_rsp_data <= 32'h05700035;
        16'h01BC : rd_rsp_data <= 32'h0154C222;
        16'h01C4 : rd_rsp_data <= 32'h00000754;
        16'h01C8 : rd_rsp_data <= 32'h78000000;
        16'h01D8 : rd_rsp_data <= 32'h07400000;
        16'h01DC : rd_rsp_data <= 32'h02180080;
        16'h01E0 : rd_rsp_data <= 32'h00162000;
        16'h01E8 : rd_rsp_data <= 32'h40000000;
        16'h0200 : rd_rsp_data <= 32'h001C1414;
        16'h0204 : rd_rsp_data <= 32'h00311414;
        16'h0208 : rd_rsp_data <= 32'h00081819;
        16'h020C : rd_rsp_data <= 32'h0024181C;
        16'h0210 : rd_rsp_data <= 32'h00211D1D;
        16'h0214 : rd_rsp_data <= 32'h00100C0C;
        16'h0218 : rd_rsp_data <= 32'h001D181C;
        16'h021C : rd_rsp_data <= 32'h000C1418;
        16'h0280 : rd_rsp_data <= 32'h10C68000;
        16'h0284 : rd_rsp_data <= 32'hF0F87843;
        16'h0288 : rd_rsp_data <= 32'hFC212480;
        16'h028C : rd_rsp_data <= 32'h0053C001;
        16'h0290 : rd_rsp_data <= 32'h4F1E1000;
        16'h0294 : rd_rsp_data <= 32'h00063C21;
        16'h0298 : rd_rsp_data <= 32'h4FE00000;
        16'h029C : rd_rsp_data <= 32'h0A025B81;
        16'h02A0 : rd_rsp_data <= 32'h9FF0577E;
        16'h02A4 : rd_rsp_data <= 32'h1C210FBE;
        16'h02A8 : rd_rsp_data <= 32'h98C011DF;
        16'h02AC : rd_rsp_data <= 32'hA8000000;
        16'h02B0 : rd_rsp_data <= 32'h045E4904;
        16'h02B4 : rd_rsp_data <= 32'h061C003B;
        16'h02B8 : rd_rsp_data <= 32'h8820E21F;
        16'h02BC : rd_rsp_data <= 32'h58155D63;
        16'h02C8 : rd_rsp_data <= 32'h30000000;
        16'h02D4 : rd_rsp_data <= 32'h01041041;
        16'h02D8 : rd_rsp_data <= 32'h08208080;
        16'h02DC : rd_rsp_data <= 32'h1E560820;
        16'h02E0 : rd_rsp_data <= 32'h806D4D93;
        16'h02E4 : rd_rsp_data <= 32'h68646467;
        16'h02E8 : rd_rsp_data <= 32'h80525A56;
        16'h02EC : rd_rsp_data <= 32'h80808080;
        16'h02F0 : rd_rsp_data <= 32'h80808080;
        16'h02F4 : rd_rsp_data <= 32'h01429339;
        16'h02F8 : rd_rsp_data <= 32'h01020FFF;
        16'h02FC : rd_rsp_data <= 32'h01020FFF;
        16'h0300 : rd_rsp_data <= 32'h01020FFF;
        16'h0308 : rd_rsp_data <= 32'h001F13AB;
        16'h030C : rd_rsp_data <= 32'h00FFFFFF;
        16'h0310 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0314 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0320 : rd_rsp_data <= 32'h0001A000;
        16'h0328 : rd_rsp_data <= 32'h03800000;
        16'h032C : rd_rsp_data <= 32'h076889AF;
        16'h033C : rd_rsp_data <= 32'h023600E3;
        16'h0340 : rd_rsp_data <= 32'h0006087E;
        16'h0348 : rd_rsp_data <= 32'h80100010;
        16'h034C : rd_rsp_data <= 32'h99999999;
        16'h0350 : rd_rsp_data <= 32'h21084290;
        16'h0354 : rd_rsp_data <= 32'h210842D0;
        16'h0358 : rd_rsp_data <= 32'h21084230;
        16'h035C : rd_rsp_data <= 32'h210841F0;
        16'h0360 : rd_rsp_data <= 32'h21084270;
        16'h0364 : rd_rsp_data <= 32'h21084250;
        16'h0368 : rd_rsp_data <= 32'h21084250;
        16'h036C : rd_rsp_data <= 32'h21084250;
        16'h0370 : rd_rsp_data <= 32'h21084210;
        16'h0374 : rd_rsp_data <= 32'h21084210;
        16'h0378 : rd_rsp_data <= 32'h00084210;
        16'h037C : rd_rsp_data <= 32'h00077054;
        16'h0380 : rd_rsp_data <= 32'h08400000;
        16'h0398 : rd_rsp_data <= 32'h808CF60A;
        16'h039C : rd_rsp_data <= 32'h00000016;
        16'h03A0 : rd_rsp_data <= 32'h00019400;
        16'h03AC : rd_rsp_data <= 32'h03260244;
        16'h03B0 : rd_rsp_data <= 32'h12481000;
        16'h03B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h03B8 : rd_rsp_data <= 32'h05800035;
        16'h03BC : rd_rsp_data <= 32'h0154C222;
        16'h03C4 : rd_rsp_data <= 32'h0000076E;
        16'h03C8 : rd_rsp_data <= 32'h78000000;
        16'h03D8 : rd_rsp_data <= 32'h07400000;
        16'h03DC : rd_rsp_data <= 32'h02180080;
        16'h03E0 : rd_rsp_data <= 32'h00162000;
        16'h03E8 : rd_rsp_data <= 32'h40000000;
        16'h0400 : rd_rsp_data <= 32'h00102529;
        16'h0404 : rd_rsp_data <= 32'h0025100C;
        16'h0408 : rd_rsp_data <= 32'h002D1C15;
        16'h040C : rd_rsp_data <= 32'h00252929;
        16'h0410 : rd_rsp_data <= 32'h001D1D14;
        16'h0414 : rd_rsp_data <= 32'h003A1810;
        16'h0418 : rd_rsp_data <= 32'h001C251D;
        16'h041C : rd_rsp_data <= 32'h00201C19;
        16'h0480 : rd_rsp_data <= 32'h10C68000;
        16'h0484 : rd_rsp_data <= 32'hF0F87843;
        16'h0488 : rd_rsp_data <= 32'hFC212480;
        16'h048C : rd_rsp_data <= 32'h005B0001;
        16'h0490 : rd_rsp_data <= 32'h4F9E1000;
        16'h0494 : rd_rsp_data <= 32'h00063C21;
        16'h0498 : rd_rsp_data <= 32'h4FE00000;
        16'h049C : rd_rsp_data <= 32'h0A025B81;
        16'h04A0 : rd_rsp_data <= 32'h9FF057FE;
        16'h04A4 : rd_rsp_data <= 32'h04210FBF;
        16'h04A8 : rd_rsp_data <= 32'h98C011DF;
        16'h04AC : rd_rsp_data <= 32'hA8000000;
        16'h04B0 : rd_rsp_data <= 32'h045E4904;
        16'h04B4 : rd_rsp_data <= 32'h061C003B;
        16'h04B8 : rd_rsp_data <= 32'h8820EE1F;
        16'h04BC : rd_rsp_data <= 32'h58155D63;
        16'h04C8 : rd_rsp_data <= 32'h30000000;
        16'h04D4 : rd_rsp_data <= 32'h01041041;
        16'h04D8 : rd_rsp_data <= 32'h08208080;
        16'h04DC : rd_rsp_data <= 32'h1E560820;
        16'h04E0 : rd_rsp_data <= 32'h80684E8B;
        16'h04E4 : rd_rsp_data <= 32'h6C666C5C;
        16'h04E8 : rd_rsp_data <= 32'h80616A52;
        16'h04EC : rd_rsp_data <= 32'h80808080;
        16'h04F0 : rd_rsp_data <= 32'h80808080;
        16'h04F4 : rd_rsp_data <= 32'h0142C3E7;
        16'h04F8 : rd_rsp_data <= 32'h01020FFF;
        16'h04FC : rd_rsp_data <= 32'h01020FFF;
        16'h0500 : rd_rsp_data <= 32'h01020FFF;
        16'h0508 : rd_rsp_data <= 32'h002113B7;
        16'h050C : rd_rsp_data <= 32'h00FFFFFF;
        16'h0510 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0514 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0528 : rd_rsp_data <= 32'h03800000;
        16'h052C : rd_rsp_data <= 32'h06458BBC;
        16'h053C : rd_rsp_data <= 32'h023404E3;
        16'h0540 : rd_rsp_data <= 32'h0006087E;
        16'h0548 : rd_rsp_data <= 32'h80100010;
        16'h054C : rd_rsp_data <= 32'h99999999;
        16'h0550 : rd_rsp_data <= 32'h210841D0;
        16'h0554 : rd_rsp_data <= 32'h21084210;
        16'h0558 : rd_rsp_data <= 32'h21084210;
        16'h055C : rd_rsp_data <= 32'h21084230;
        16'h0560 : rd_rsp_data <= 32'h210842D0;
        16'h0564 : rd_rsp_data <= 32'h210841F0;
        16'h0568 : rd_rsp_data <= 32'h210841F0;
        16'h056C : rd_rsp_data <= 32'h21084210;
        16'h0570 : rd_rsp_data <= 32'h21084210;
        16'h0574 : rd_rsp_data <= 32'h21084210;
        16'h0578 : rd_rsp_data <= 32'h00084210;
        16'h057C : rd_rsp_data <= 32'h00077054;
        16'h0580 : rd_rsp_data <= 32'h08400000;
        16'h0598 : rd_rsp_data <= 32'h808CF60A;
        16'h059C : rd_rsp_data <= 32'h00000016;
        16'h05A0 : rd_rsp_data <= 32'h00019400;
        16'h05AC : rd_rsp_data <= 32'h03260244;
        16'h05B0 : rd_rsp_data <= 32'h12481000;
        16'h05B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h05B8 : rd_rsp_data <= 32'h05800035;
        16'h05BC : rd_rsp_data <= 32'h0154C222;
        16'h05C4 : rd_rsp_data <= 32'h000007EC;
        16'h05C8 : rd_rsp_data <= 32'h78000000;
        16'h05D8 : rd_rsp_data <= 32'h07400000;
        16'h05DC : rd_rsp_data <= 32'h02180080;
        16'h05E0 : rd_rsp_data <= 32'h00162000;
        16'h05E8 : rd_rsp_data <= 32'h40000000;
        16'h0600 : rd_rsp_data <= 32'h0010191C;
        16'h0604 : rd_rsp_data <= 32'h0024191C;
        16'h0608 : rd_rsp_data <= 32'h00181410;
        16'h060C : rd_rsp_data <= 32'h00291818;
        16'h0610 : rd_rsp_data <= 32'h002E0810;
        16'h0614 : rd_rsp_data <= 32'h00210C10;
        16'h0618 : rd_rsp_data <= 32'h00140C14;
        16'h061C : rd_rsp_data <= 32'h00101014;
        16'h0680 : rd_rsp_data <= 32'h10C68000;
        16'h0684 : rd_rsp_data <= 32'hF0F87843;
        16'h0688 : rd_rsp_data <= 32'hFC212480;
        16'h068C : rd_rsp_data <= 32'h005AC001;
        16'h0690 : rd_rsp_data <= 32'h4F1E1000;
        16'h0694 : rd_rsp_data <= 32'h00063C21;
        16'h0698 : rd_rsp_data <= 32'h4EE00000;
        16'h069C : rd_rsp_data <= 32'h0A025B81;
        16'h06A0 : rd_rsp_data <= 32'h9FF057BC;
        16'h06A4 : rd_rsp_data <= 32'h84210FFE;
        16'h06A8 : rd_rsp_data <= 32'h98C011DF;
        16'h06AC : rd_rsp_data <= 32'hA8000000;
        16'h06B0 : rd_rsp_data <= 32'h045E4904;
        16'h06B4 : rd_rsp_data <= 32'h061C003B;
        16'h06B8 : rd_rsp_data <= 32'h8820EE1F;
        16'h06BC : rd_rsp_data <= 32'h58155D63;
        16'h06C8 : rd_rsp_data <= 32'h30000000;
        16'h06D4 : rd_rsp_data <= 32'h01041041;
        16'h06D8 : rd_rsp_data <= 32'h08208080;
        16'h06DC : rd_rsp_data <= 32'h1E560820;
        16'h06E0 : rd_rsp_data <= 32'h806C6A83;
        16'h06E4 : rd_rsp_data <= 32'h64746E6D;
        16'h06E8 : rd_rsp_data <= 32'h80625A50;
        16'h06EC : rd_rsp_data <= 32'h80808080;
        16'h06F0 : rd_rsp_data <= 32'h80808080;
        16'h06F4 : rd_rsp_data <= 32'h014AA333;
        16'h06F8 : rd_rsp_data <= 32'h01020FFF;
        16'h06FC : rd_rsp_data <= 32'h01020FFF;
        16'h0700 : rd_rsp_data <= 32'h01020FFF;
        16'h0708 : rd_rsp_data <= 32'h001E939D;
        16'h070C : rd_rsp_data <= 32'h00FFFFFF;
        16'h0710 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0714 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0728 : rd_rsp_data <= 32'h03800000;
        16'h072C : rd_rsp_data <= 32'h066889AF;
        16'h073C : rd_rsp_data <= 32'h023600E3;
        16'h0740 : rd_rsp_data <= 32'h0006087E;
        16'h0748 : rd_rsp_data <= 32'h80100010;
        16'h074C : rd_rsp_data <= 32'h99999999;
        16'h0750 : rd_rsp_data <= 32'h21084250;
        16'h0754 : rd_rsp_data <= 32'h21084250;
        16'h0758 : rd_rsp_data <= 32'h21084230;
        16'h075C : rd_rsp_data <= 32'h210841F0;
        16'h0760 : rd_rsp_data <= 32'h21084270;
        16'h0764 : rd_rsp_data <= 32'h21084270;
        16'h0768 : rd_rsp_data <= 32'h21084230;
        16'h076C : rd_rsp_data <= 32'h21084270;
        16'h0770 : rd_rsp_data <= 32'h21084210;
        16'h0774 : rd_rsp_data <= 32'h21084210;
        16'h0778 : rd_rsp_data <= 32'h00084210;
        16'h077C : rd_rsp_data <= 32'h00077054;
        16'h0780 : rd_rsp_data <= 32'h08400000;
        16'h0798 : rd_rsp_data <= 32'h808CF60A;
        16'h079C : rd_rsp_data <= 32'h00000016;
        16'h07A0 : rd_rsp_data <= 32'h00019400;
        16'h07AC : rd_rsp_data <= 32'h03260244;
        16'h07B0 : rd_rsp_data <= 32'h12481000;
        16'h07B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h07B8 : rd_rsp_data <= 32'h05800035;
        16'h07BC : rd_rsp_data <= 32'h0154C222;
        16'h07C4 : rd_rsp_data <= 32'h00000016;
        16'h07C8 : rd_rsp_data <= 32'h78000000;
        16'h07D8 : rd_rsp_data <= 32'h07400000;
        16'h07DC : rd_rsp_data <= 32'h02180080;
        16'h07E0 : rd_rsp_data <= 32'h00162000;
        16'h07E8 : rd_rsp_data <= 32'h40000000;
        16'h0800 : rd_rsp_data <= 32'h0014100C;
        16'h0804 : rd_rsp_data <= 32'h00101D10;
        16'h0808 : rd_rsp_data <= 32'h00291414;
        16'h080C : rd_rsp_data <= 32'h00291008;
        16'h0810 : rd_rsp_data <= 32'h00251004;
        16'h0814 : rd_rsp_data <= 32'h0028140C;
        16'h0818 : rd_rsp_data <= 32'h00101814;
        16'h081C : rd_rsp_data <= 32'h001C2519;
        16'h0880 : rd_rsp_data <= 32'h10C68000;
        16'h0884 : rd_rsp_data <= 32'hF0F87843;
        16'h0888 : rd_rsp_data <= 32'hFC212480;
        16'h088C : rd_rsp_data <= 32'h005A0001;
        16'h0890 : rd_rsp_data <= 32'h4F1E1000;
        16'h0894 : rd_rsp_data <= 32'h00063C21;
        16'h0898 : rd_rsp_data <= 32'h4EE00000;
        16'h089C : rd_rsp_data <= 32'h0A025B81;
        16'h08A0 : rd_rsp_data <= 32'h9FF057BE;
        16'h08A4 : rd_rsp_data <= 32'hAC210FBF;
        16'h08A8 : rd_rsp_data <= 32'h98C011DF;
        16'h08AC : rd_rsp_data <= 32'hA8000000;
        16'h08B0 : rd_rsp_data <= 32'h045E4904;
        16'h08B4 : rd_rsp_data <= 32'h061C003B;
        16'h08B8 : rd_rsp_data <= 32'h8820F21F;
        16'h08BC : rd_rsp_data <= 32'h58155D63;
        16'h08C8 : rd_rsp_data <= 32'h30000000;
        16'h08D4 : rd_rsp_data <= 32'h01041041;
        16'h08D8 : rd_rsp_data <= 32'h08208080;
        16'h08DC : rd_rsp_data <= 32'h1E560820;
        16'h08E0 : rd_rsp_data <= 32'h804A5684;
        16'h08E4 : rd_rsp_data <= 32'h4B4A585E;
        16'h08E8 : rd_rsp_data <= 32'h80504F4A;
        16'h08EC : rd_rsp_data <= 32'h80808080;
        16'h08F0 : rd_rsp_data <= 32'h80808080;
        16'h08F4 : rd_rsp_data <= 32'h0162E37D;
        16'h08F8 : rd_rsp_data <= 32'h01020FFF;
        16'h08FC : rd_rsp_data <= 32'h01020FFF;
        16'h0900 : rd_rsp_data <= 32'h01020FFF;
        16'h0908 : rd_rsp_data <= 32'h001C5371;
        16'h090C : rd_rsp_data <= 32'h00FFFFFF;
        16'h0910 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0914 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0928 : rd_rsp_data <= 32'h03800000;
        16'h092C : rd_rsp_data <= 32'h0744397E;
        16'h093C : rd_rsp_data <= 32'h023C04E0;
        16'h0940 : rd_rsp_data <= 32'h0006087E;
        16'h0948 : rd_rsp_data <= 32'h80100010;
        16'h094C : rd_rsp_data <= 32'h99999999;
        16'h0950 : rd_rsp_data <= 32'h21084290;
        16'h0954 : rd_rsp_data <= 32'h210842F0;
        16'h0958 : rd_rsp_data <= 32'h21084230;
        16'h095C : rd_rsp_data <= 32'h21084230;
        16'h0960 : rd_rsp_data <= 32'h210841F0;
        16'h0964 : rd_rsp_data <= 32'h21084230;
        16'h0968 : rd_rsp_data <= 32'h21084250;
        16'h096C : rd_rsp_data <= 32'h21084250;
        16'h0970 : rd_rsp_data <= 32'h21084210;
        16'h0974 : rd_rsp_data <= 32'h21084210;
        16'h0978 : rd_rsp_data <= 32'h00084210;
        16'h097C : rd_rsp_data <= 32'h00077054;
        16'h0980 : rd_rsp_data <= 32'h08400000;
        16'h0998 : rd_rsp_data <= 32'h808CF60A;
        16'h099C : rd_rsp_data <= 32'h00000016;
        16'h09A0 : rd_rsp_data <= 32'h00019400;
        16'h09AC : rd_rsp_data <= 32'h03260244;
        16'h09B0 : rd_rsp_data <= 32'h12481000;
        16'h09B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h09B8 : rd_rsp_data <= 32'h05800035;
        16'h09BC : rd_rsp_data <= 32'h0154C222;
        16'h09C4 : rd_rsp_data <= 32'h000006FE;
        16'h09C8 : rd_rsp_data <= 32'h78000000;
        16'h09D8 : rd_rsp_data <= 32'h07400000;
        16'h09DC : rd_rsp_data <= 32'h02180080;
        16'h09E0 : rd_rsp_data <= 32'h00162000;
        16'h09E8 : rd_rsp_data <= 32'h40000000;
        16'h0A00 : rd_rsp_data <= 32'h0028140C;
        16'h0A04 : rd_rsp_data <= 32'h00311410;
        16'h0A08 : rd_rsp_data <= 32'h00141814;
        16'h0A0C : rd_rsp_data <= 32'h00291814;
        16'h0A10 : rd_rsp_data <= 32'h00101810;
        16'h0A14 : rd_rsp_data <= 32'h00201010;
        16'h0A18 : rd_rsp_data <= 32'h00241818;
        16'h0A1C : rd_rsp_data <= 32'h00181410;
        16'h0A80 : rd_rsp_data <= 32'h10C68000;
        16'h0A84 : rd_rsp_data <= 32'hF0783801;
        16'h0A88 : rd_rsp_data <= 32'hFC212480;
        16'h0A8C : rd_rsp_data <= 32'h00578001;
        16'h0A90 : rd_rsp_data <= 32'h4F1E1000;
        16'h0A94 : rd_rsp_data <= 32'h00063C21;
        16'h0A98 : rd_rsp_data <= 32'h4FE00000;
        16'h0A9C : rd_rsp_data <= 32'h0A025B81;
        16'h0AA0 : rd_rsp_data <= 32'h9FF05778;
        16'h0AA4 : rd_rsp_data <= 32'hE4210FFA;
        16'h0AA8 : rd_rsp_data <= 32'h98C011DF;
        16'h0AAC : rd_rsp_data <= 32'hA8000000;
        16'h0AB0 : rd_rsp_data <= 32'h045E4904;
        16'h0AB4 : rd_rsp_data <= 32'h061C003B;
        16'h0AB8 : rd_rsp_data <= 32'h8820F21F;
        16'h0ABC : rd_rsp_data <= 32'h58155D63;
        16'h0AC8 : rd_rsp_data <= 32'h30000000;
        16'h0AD4 : rd_rsp_data <= 32'h01041041;
        16'h0AD8 : rd_rsp_data <= 32'h08208080;
        16'h0ADC : rd_rsp_data <= 32'h1E560820;
        16'h0AE0 : rd_rsp_data <= 32'h80785793;
        16'h0AE4 : rd_rsp_data <= 32'h69787369;
        16'h0AE8 : rd_rsp_data <= 32'h807C6464;
        16'h0AEC : rd_rsp_data <= 32'h80808080;
        16'h0AF0 : rd_rsp_data <= 32'h80808080;
        16'h0AF4 : rd_rsp_data <= 32'h0152A2AF;
        16'h0AF8 : rd_rsp_data <= 32'h01020FFF;
        16'h0AFC : rd_rsp_data <= 32'h01020FFF;
        16'h0B00 : rd_rsp_data <= 32'h01020FFF;
        16'h0B08 : rd_rsp_data <= 32'h001B9367;
        16'h0B0C : rd_rsp_data <= 32'h00FFFFFF;
        16'h0B10 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0B14 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0B20 : rd_rsp_data <= 32'h0001D000;
        16'h0B28 : rd_rsp_data <= 32'h03800000;
        16'h0B2C : rd_rsp_data <= 32'h0705A9BD;
        16'h0B3C : rd_rsp_data <= 32'h023200E5;
        16'h0B40 : rd_rsp_data <= 32'h0006087E;
        16'h0B48 : rd_rsp_data <= 32'h80100010;
        16'h0B4C : rd_rsp_data <= 32'h99999999;
        16'h0B50 : rd_rsp_data <= 32'h210842D0;
        16'h0B54 : rd_rsp_data <= 32'h21084230;
        16'h0B58 : rd_rsp_data <= 32'h21084290;
        16'h0B5C : rd_rsp_data <= 32'h21084290;
        16'h0B60 : rd_rsp_data <= 32'h210842F0;
        16'h0B64 : rd_rsp_data <= 32'h21084210;
        16'h0B68 : rd_rsp_data <= 32'h21084230;
        16'h0B6C : rd_rsp_data <= 32'h21084230;
        16'h0B70 : rd_rsp_data <= 32'h21084210;
        16'h0B74 : rd_rsp_data <= 32'h21084210;
        16'h0B78 : rd_rsp_data <= 32'h00084210;
        16'h0B7C : rd_rsp_data <= 32'h00077054;
        16'h0B80 : rd_rsp_data <= 32'h08400000;
        16'h0B98 : rd_rsp_data <= 32'h808CF60A;
        16'h0B9C : rd_rsp_data <= 32'h00000016;
        16'h0BA0 : rd_rsp_data <= 32'h00019400;
        16'h0BAC : rd_rsp_data <= 32'h03260244;
        16'h0BB0 : rd_rsp_data <= 32'h12481000;
        16'h0BB4 : rd_rsp_data <= 32'h2D495C3E;
        16'h0BB8 : rd_rsp_data <= 32'h05800035;
        16'h0BBC : rd_rsp_data <= 32'h0154C222;
        16'h0BC4 : rd_rsp_data <= 32'h0000077A;
        16'h0BC8 : rd_rsp_data <= 32'h78000000;
        16'h0BD8 : rd_rsp_data <= 32'h07400000;
        16'h0BDC : rd_rsp_data <= 32'h02180080;
        16'h0BE0 : rd_rsp_data <= 32'h00162000;
        16'h0BE8 : rd_rsp_data <= 32'h40000000;
        16'h0C00 : rd_rsp_data <= 32'h00291914;
        16'h0C04 : rd_rsp_data <= 32'h0025100C;
        16'h0C08 : rd_rsp_data <= 32'h00320804;
        16'h0C0C : rd_rsp_data <= 32'h00141819;
        16'h0C10 : rd_rsp_data <= 32'h002D2115;
        16'h0C14 : rd_rsp_data <= 32'h0031100C;
        16'h0C18 : rd_rsp_data <= 32'h0010211D;
        16'h0C1C : rd_rsp_data <= 32'h00211D14;
        16'h0C80 : rd_rsp_data <= 32'h10C68000;
        16'h0C84 : rd_rsp_data <= 32'hF0F87843;
        16'h0C88 : rd_rsp_data <= 32'hFC212480;
        16'h0C8C : rd_rsp_data <= 32'h005BC001;
        16'h0C90 : rd_rsp_data <= 32'h4F9E1000;
        16'h0C94 : rd_rsp_data <= 32'h00063C21;
        16'h0C98 : rd_rsp_data <= 32'h5DE00000;
        16'h0C9C : rd_rsp_data <= 32'h0A025B81;
        16'h0CA0 : rd_rsp_data <= 32'h9FF057BE;
        16'h0CA4 : rd_rsp_data <= 32'h9C210FBF;
        16'h0CA8 : rd_rsp_data <= 32'h98C011DF;
        16'h0CAC : rd_rsp_data <= 32'hA8000000;
        16'h0CB0 : rd_rsp_data <= 32'h045E4904;
        16'h0CB4 : rd_rsp_data <= 32'h061C003B;
        16'h0CB8 : rd_rsp_data <= 32'h8820E61F;
        16'h0CBC : rd_rsp_data <= 32'h58155D63;
        16'h0CC8 : rd_rsp_data <= 32'h30000000;
        16'h0CD4 : rd_rsp_data <= 32'h01041041;
        16'h0CD8 : rd_rsp_data <= 32'h08208080;
        16'h0CDC : rd_rsp_data <= 32'h1E560820;
        16'h0CE0 : rd_rsp_data <= 32'h80785480;
        16'h0CE4 : rd_rsp_data <= 32'h7A807C70;
        16'h0CE8 : rd_rsp_data <= 32'h8072706B;
        16'h0CEC : rd_rsp_data <= 32'h80808080;
        16'h0CF0 : rd_rsp_data <= 32'h80808080;
        16'h0CF4 : rd_rsp_data <= 32'h014AC36D;
        16'h0CF8 : rd_rsp_data <= 32'h01020FFF;
        16'h0CFC : rd_rsp_data <= 32'h01020FFF;
        16'h0D00 : rd_rsp_data <= 32'h01020FFF;
        16'h0D08 : rd_rsp_data <= 32'h001D1379;
        16'h0D0C : rd_rsp_data <= 32'h00FFFFFF;
        16'h0D10 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0D14 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0D20 : rd_rsp_data <= 32'h00003000;
        16'h0D28 : rd_rsp_data <= 32'h03800000;
        16'h0D2C : rd_rsp_data <= 32'h0644397E;
        16'h0D3C : rd_rsp_data <= 32'h023C04E0;
        16'h0D40 : rd_rsp_data <= 32'h0006087E;
        16'h0D48 : rd_rsp_data <= 32'h80100010;
        16'h0D4C : rd_rsp_data <= 32'h99999999;
        16'h0D50 : rd_rsp_data <= 32'h21084230;
        16'h0D54 : rd_rsp_data <= 32'h21084210;
        16'h0D58 : rd_rsp_data <= 32'h21084210;
        16'h0D5C : rd_rsp_data <= 32'h210842D0;
        16'h0D60 : rd_rsp_data <= 32'h21084250;
        16'h0D64 : rd_rsp_data <= 32'h21084230;
        16'h0D68 : rd_rsp_data <= 32'h21084250;
        16'h0D6C : rd_rsp_data <= 32'h210841F0;
        16'h0D70 : rd_rsp_data <= 32'h21084210;
        16'h0D74 : rd_rsp_data <= 32'h21084210;
        16'h0D78 : rd_rsp_data <= 32'h00084210;
        16'h0D7C : rd_rsp_data <= 32'h00077054;
        16'h0D80 : rd_rsp_data <= 32'h08400000;
        16'h0D98 : rd_rsp_data <= 32'h808CF60A;
        16'h0D9C : rd_rsp_data <= 32'h00000012;
        16'h0DA0 : rd_rsp_data <= 32'h00019400;
        16'h0DAC : rd_rsp_data <= 32'h03260244;
        16'h0DB0 : rd_rsp_data <= 32'h12481000;
        16'h0DB4 : rd_rsp_data <= 32'h2D495C3E;
        16'h0DB8 : rd_rsp_data <= 32'h05800035;
        16'h0DBC : rd_rsp_data <= 32'h0154C222;
        16'h0DC4 : rd_rsp_data <= 32'h000006EE;
        16'h0DC8 : rd_rsp_data <= 32'h78000000;
        16'h0DD8 : rd_rsp_data <= 32'h07400000;
        16'h0DDC : rd_rsp_data <= 32'h02180080;
        16'h0DE0 : rd_rsp_data <= 32'h00122000;
        16'h0DE8 : rd_rsp_data <= 32'h40000000;
        16'h0E00 : rd_rsp_data <= 32'h003A1819;
        16'h0E04 : rd_rsp_data <= 32'h001C100C;
        16'h0E08 : rd_rsp_data <= 32'h00181018;
        16'h0E0C : rd_rsp_data <= 32'h00311015;
        16'h0E10 : rd_rsp_data <= 32'h00290C15;
        16'h0E14 : rd_rsp_data <= 32'h000C1010;
        16'h0E18 : rd_rsp_data <= 32'h00210C15;
        16'h0E1C : rd_rsp_data <= 32'h00201419;
        16'h0E80 : rd_rsp_data <= 32'h10C68000;
        16'h0E84 : rd_rsp_data <= 32'hF0783801;
        16'h0E88 : rd_rsp_data <= 32'hFC212480;
        16'h0E8C : rd_rsp_data <= 32'h00580001;
        16'h0E90 : rd_rsp_data <= 32'h4D1E1000;
        16'h0E94 : rd_rsp_data <= 32'h00063C21;
        16'h0E98 : rd_rsp_data <= 32'h4FE00000;
        16'h0E9C : rd_rsp_data <= 32'h0A025B81;
        16'h0EA0 : rd_rsp_data <= 32'h9FF057F8;
        16'h0EA4 : rd_rsp_data <= 32'h8C210FFE;
        16'h0EA8 : rd_rsp_data <= 32'h98C011DF;
        16'h0EAC : rd_rsp_data <= 32'hA8000000;
        16'h0EB0 : rd_rsp_data <= 32'h045E4904;
        16'h0EB4 : rd_rsp_data <= 32'h061C003B;
        16'h0EB8 : rd_rsp_data <= 32'h8820EE1F;
        16'h0EBC : rd_rsp_data <= 32'h58155D63;
        16'h0EC8 : rd_rsp_data <= 32'h30000000;
        16'h0ED4 : rd_rsp_data <= 32'h01041041;
        16'h0ED8 : rd_rsp_data <= 32'h08208080;
        16'h0EDC : rd_rsp_data <= 32'h1E560820;
        16'h0EE0 : rd_rsp_data <= 32'h806C528B;
        16'h0EE4 : rd_rsp_data <= 32'h68586C5C;
        16'h0EE8 : rd_rsp_data <= 32'h80706065;
        16'h0EEC : rd_rsp_data <= 32'h80808080;
        16'h0EF0 : rd_rsp_data <= 32'h80808080;
        16'h0EF4 : rd_rsp_data <= 32'h015282A9;
        16'h0EF8 : rd_rsp_data <= 32'h01020FFF;
        16'h0EFC : rd_rsp_data <= 32'h01020FFF;
        16'h0F00 : rd_rsp_data <= 32'h01020FFF;
        16'h0F08 : rd_rsp_data <= 32'h001C1373;
        16'h0F0C : rd_rsp_data <= 32'h00FFFFFF;
        16'h0F10 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0F14 : rd_rsp_data <= 32'h00FFFFFF;
        16'h0F20 : rd_rsp_data <= 32'h0001D000;
        16'h0F28 : rd_rsp_data <= 32'h03800000;
        16'h0F2C : rd_rsp_data <= 32'h0605A9BD;
        16'h0F3C : rd_rsp_data <= 32'h023200E5;
        16'h0F40 : rd_rsp_data <= 32'h0006087E;
        16'h0F48 : rd_rsp_data <= 32'h80100010;
        16'h0F4C : rd_rsp_data <= 32'h99999999;
        16'h0F50 : rd_rsp_data <= 32'h21084330;
        16'h0F54 : rd_rsp_data <= 32'h21084290;
        16'h0F58 : rd_rsp_data <= 32'h21084270;
        16'h0F5C : rd_rsp_data <= 32'h21084210;
        16'h0F60 : rd_rsp_data <= 32'h21084270;
        16'h0F64 : rd_rsp_data <= 32'h21084210;
        16'h0F68 : rd_rsp_data <= 32'h21084310;
        16'h0F6C : rd_rsp_data <= 32'h21084250;
        16'h0F70 : rd_rsp_data <= 32'h21084210;
        16'h0F74 : rd_rsp_data <= 32'h21084210;
        16'h0F78 : rd_rsp_data <= 32'h00084210;
        16'h0F7C : rd_rsp_data <= 32'h00077054;
        16'h0F80 : rd_rsp_data <= 32'h08400000;
        16'h0F98 : rd_rsp_data <= 32'h808CF60A;
        16'h0F9C : rd_rsp_data <= 32'h00000016;
        16'h0FA0 : rd_rsp_data <= 32'h00019400;
        16'h0FAC : rd_rsp_data <= 32'h03260244;
        16'h0FB0 : rd_rsp_data <= 32'h12481000;
        16'h0FB4 : rd_rsp_data <= 32'h2D495C3E;
        16'h0FB8 : rd_rsp_data <= 32'h05800035;
        16'h0FBC : rd_rsp_data <= 32'h0154C222;
        16'h0FC4 : rd_rsp_data <= 32'h0000031C;
        16'h0FC8 : rd_rsp_data <= 32'h7F000000;
        16'h0FD8 : rd_rsp_data <= 32'h07400000;
        16'h0FDC : rd_rsp_data <= 32'h02180080;
        16'h0FE0 : rd_rsp_data <= 32'h00162000;
        16'h0FE8 : rd_rsp_data <= 32'h40000000;
        16'h1000 : rd_rsp_data <= 32'h00421D18;
        16'h1004 : rd_rsp_data <= 32'h002D0C0C;
        16'h1008 : rd_rsp_data <= 32'h003A1010;
        16'h100C : rd_rsp_data <= 32'h0025080C;
        16'h1010 : rd_rsp_data <= 32'h00351818;
        16'h1014 : rd_rsp_data <= 32'h00361818;
        16'h1018 : rd_rsp_data <= 32'h00182929;
        16'h101C : rd_rsp_data <= 32'h00351010;
        16'h1080 : rd_rsp_data <= 32'h10C68000;
        16'h1084 : rd_rsp_data <= 32'hF0F87843;
        16'h1088 : rd_rsp_data <= 32'hFC212480;
        16'h108C : rd_rsp_data <= 32'h005AC001;
        16'h1090 : rd_rsp_data <= 32'h4F9E1000;
        16'h1094 : rd_rsp_data <= 32'h00063C21;
        16'h1098 : rd_rsp_data <= 32'h4EE00000;
        16'h109C : rd_rsp_data <= 32'h0A025B81;
        16'h10A0 : rd_rsp_data <= 32'h9FF054FE;
        16'h10A4 : rd_rsp_data <= 32'h54210F76;
        16'h10A8 : rd_rsp_data <= 32'h98C011DF;
        16'h10AC : rd_rsp_data <= 32'hA8000000;
        16'h10B0 : rd_rsp_data <= 32'h045E4904;
        16'h10B4 : rd_rsp_data <= 32'h061C003B;
        16'h10B8 : rd_rsp_data <= 32'h8820EE1F;
        16'h10BC : rd_rsp_data <= 32'h58155D63;
        16'h10C8 : rd_rsp_data <= 32'h30000000;
        16'h10D4 : rd_rsp_data <= 32'h01041041;
        16'h10D8 : rd_rsp_data <= 32'h08208080;
        16'h10DC : rd_rsp_data <= 32'h1E560820;
        16'h10E0 : rd_rsp_data <= 32'h8062788B;
        16'h10E4 : rd_rsp_data <= 32'h745A6E72;
        16'h10E8 : rd_rsp_data <= 32'h80635C5C;
        16'h10EC : rd_rsp_data <= 32'h80808080;
        16'h10F0 : rd_rsp_data <= 32'h80808080;
        16'h10F4 : rd_rsp_data <= 32'h015AB343;
        16'h10F8 : rd_rsp_data <= 32'h01020FFF;
        16'h10FC : rd_rsp_data <= 32'h01020FFF;
        16'h1100 : rd_rsp_data <= 32'h01020FFF;
        16'h1108 : rd_rsp_data <= 32'h001D537F;
        16'h110C : rd_rsp_data <= 32'h00FFFFFF;
        16'h1110 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1114 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1128 : rd_rsp_data <= 32'h03800000;
        16'h112C : rd_rsp_data <= 32'h060D19EE;
        16'h113C : rd_rsp_data <= 32'h023000E5;
        16'h1140 : rd_rsp_data <= 32'h0006087E;
        16'h1148 : rd_rsp_data <= 32'h80100010;
        16'h114C : rd_rsp_data <= 32'h99999999;
        16'h1150 : rd_rsp_data <= 32'h210842F0;
        16'h1154 : rd_rsp_data <= 32'h210842F0;
        16'h1158 : rd_rsp_data <= 32'h210842B0;
        16'h115C : rd_rsp_data <= 32'h210842B0;
        16'h1160 : rd_rsp_data <= 32'h21084190;
        16'h1164 : rd_rsp_data <= 32'h210842B0;
        16'h1168 : rd_rsp_data <= 32'h21084270;
        16'h116C : rd_rsp_data <= 32'h21084210;
        16'h1170 : rd_rsp_data <= 32'h21084210;
        16'h1174 : rd_rsp_data <= 32'h21084210;
        16'h1178 : rd_rsp_data <= 32'h00084210;
        16'h117C : rd_rsp_data <= 32'h00077054;
        16'h1180 : rd_rsp_data <= 32'h08400000;
        16'h1198 : rd_rsp_data <= 32'h808CF60A;
        16'h119C : rd_rsp_data <= 32'h00000014;
        16'h11A0 : rd_rsp_data <= 32'h00019400;
        16'h11AC : rd_rsp_data <= 32'h03260244;
        16'h11B0 : rd_rsp_data <= 32'h12481000;
        16'h11B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h11B8 : rd_rsp_data <= 32'h05800035;
        16'h11BC : rd_rsp_data <= 32'h0154C222;
        16'h11C4 : rd_rsp_data <= 32'h000003F4;
        16'h11C8 : rd_rsp_data <= 32'h78000000;
        16'h11D8 : rd_rsp_data <= 32'h07400000;
        16'h11DC : rd_rsp_data <= 32'h02180080;
        16'h11E0 : rd_rsp_data <= 32'h00142000;
        16'h11E8 : rd_rsp_data <= 32'h40000000;
        16'h1200 : rd_rsp_data <= 32'h00322114;
        16'h1204 : rd_rsp_data <= 32'h00181810;
        16'h1208 : rd_rsp_data <= 32'h003E1C10;
        16'h120C : rd_rsp_data <= 32'h001C1818;
        16'h1210 : rd_rsp_data <= 32'h00101C18;
        16'h1214 : rd_rsp_data <= 32'h00281910;
        16'h1218 : rd_rsp_data <= 32'h00251414;
        16'h121C : rd_rsp_data <= 32'h00291008;
        16'h1280 : rd_rsp_data <= 32'h10C68000;
        16'h1284 : rd_rsp_data <= 32'hF0783801;
        16'h1288 : rd_rsp_data <= 32'hFC212480;
        16'h128C : rd_rsp_data <= 32'h005DC001;
        16'h1290 : rd_rsp_data <= 32'h4E9E1000;
        16'h1294 : rd_rsp_data <= 32'h00063C21;
        16'h1298 : rd_rsp_data <= 32'h5DE00000;
        16'h129C : rd_rsp_data <= 32'h0A025B81;
        16'h12A0 : rd_rsp_data <= 32'h9FF056FE;
        16'h12A4 : rd_rsp_data <= 32'hAC210F9E;
        16'h12A8 : rd_rsp_data <= 32'h98C011DF;
        16'h12AC : rd_rsp_data <= 32'hA8000000;
        16'h12B0 : rd_rsp_data <= 32'h045E4904;
        16'h12B4 : rd_rsp_data <= 32'h061C003B;
        16'h12B8 : rd_rsp_data <= 32'h8820EE1F;
        16'h12BC : rd_rsp_data <= 32'h58155D63;
        16'h12C8 : rd_rsp_data <= 32'h30000000;
        16'h12D4 : rd_rsp_data <= 32'h01041041;
        16'h12D8 : rd_rsp_data <= 32'h08208080;
        16'h12DC : rd_rsp_data <= 32'h1E560820;
        16'h12E0 : rd_rsp_data <= 32'h80624C8B;
        16'h12E4 : rd_rsp_data <= 32'h6E685F5C;
        16'h12E8 : rd_rsp_data <= 32'h80706966;
        16'h12EC : rd_rsp_data <= 32'h80808080;
        16'h12F0 : rd_rsp_data <= 32'h80808080;
        16'h12F4 : rd_rsp_data <= 32'h0162D2A1;
        16'h12F8 : rd_rsp_data <= 32'h01020FFF;
        16'h12FC : rd_rsp_data <= 32'h01020FFF;
        16'h1300 : rd_rsp_data <= 32'h01020FFF;
        16'h1308 : rd_rsp_data <= 32'h001C1363;
        16'h130C : rd_rsp_data <= 32'h00FFFFFF;
        16'h1310 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1314 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1320 : rd_rsp_data <= 32'h00006000;
        16'h1328 : rd_rsp_data <= 32'h03800000;
        16'h132C : rd_rsp_data <= 32'h064C1D7C;
        16'h133C : rd_rsp_data <= 32'h024604DC;
        16'h1340 : rd_rsp_data <= 32'h0006087E;
        16'h1348 : rd_rsp_data <= 32'h80100010;
        16'h134C : rd_rsp_data <= 32'h99999999;
        16'h1350 : rd_rsp_data <= 32'h21084210;
        16'h1354 : rd_rsp_data <= 32'h210842B0;
        16'h1358 : rd_rsp_data <= 32'h21084250;
        16'h135C : rd_rsp_data <= 32'h21084310;
        16'h1360 : rd_rsp_data <= 32'h21084210;
        16'h1364 : rd_rsp_data <= 32'h21084330;
        16'h1368 : rd_rsp_data <= 32'h21084270;
        16'h136C : rd_rsp_data <= 32'h21084230;
        16'h1370 : rd_rsp_data <= 32'h21084210;
        16'h1374 : rd_rsp_data <= 32'h21084210;
        16'h1378 : rd_rsp_data <= 32'h00084210;
        16'h137C : rd_rsp_data <= 32'h00077054;
        16'h1380 : rd_rsp_data <= 32'h08400000;
        16'h1398 : rd_rsp_data <= 32'h808CF60A;
        16'h139C : rd_rsp_data <= 32'h00000015;
        16'h13A0 : rd_rsp_data <= 32'h00019400;
        16'h13AC : rd_rsp_data <= 32'h03260244;
        16'h13B0 : rd_rsp_data <= 32'h12481000;
        16'h13B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h13B8 : rd_rsp_data <= 32'h05800035;
        16'h13BC : rd_rsp_data <= 32'h0154C222;
        16'h13C4 : rd_rsp_data <= 32'h000007A2;
        16'h13C8 : rd_rsp_data <= 32'h7F000000;
        16'h13D8 : rd_rsp_data <= 32'h07400000;
        16'h13DC : rd_rsp_data <= 32'h02180080;
        16'h13E0 : rd_rsp_data <= 32'h00152000;
        16'h13E8 : rd_rsp_data <= 32'h40000000;
        16'h1400 : rd_rsp_data <= 32'h00311921;
        16'h1404 : rd_rsp_data <= 32'h003E0810;
        16'h1408 : rd_rsp_data <= 32'h002D0C04;
        16'h140C : rd_rsp_data <= 32'h001C0C10;
        16'h1410 : rd_rsp_data <= 32'h002D101D;
        16'h1414 : rd_rsp_data <= 32'h0020181D;
        16'h1418 : rd_rsp_data <= 32'h0029252E;
        16'h141C : rd_rsp_data <= 32'h00182125;
        16'h1480 : rd_rsp_data <= 32'h10C68000;
        16'h1484 : rd_rsp_data <= 32'hF0F87843;
        16'h1488 : rd_rsp_data <= 32'hFC212480;
        16'h148C : rd_rsp_data <= 32'h005B4001;
        16'h1490 : rd_rsp_data <= 32'h4F9E1000;
        16'h1494 : rd_rsp_data <= 32'h00063C21;
        16'h1498 : rd_rsp_data <= 32'h5DE00000;
        16'h149C : rd_rsp_data <= 32'h0A025B81;
        16'h14A0 : rd_rsp_data <= 32'h9FF057FE;
        16'h14A4 : rd_rsp_data <= 32'h24210FFD;
        16'h14A8 : rd_rsp_data <= 32'h98C011DF;
        16'h14AC : rd_rsp_data <= 32'hA8000000;
        16'h14B0 : rd_rsp_data <= 32'h045E4904;
        16'h14B4 : rd_rsp_data <= 32'h061C003B;
        16'h14B8 : rd_rsp_data <= 32'h8820F21F;
        16'h14BC : rd_rsp_data <= 32'h58155D63;
        16'h14C8 : rd_rsp_data <= 32'h30000000;
        16'h14D4 : rd_rsp_data <= 32'h01041041;
        16'h14D8 : rd_rsp_data <= 32'h08208080;
        16'h14DC : rd_rsp_data <= 32'h1E560820;
        16'h14E0 : rd_rsp_data <= 32'h805C5E9B;
        16'h14E4 : rd_rsp_data <= 32'h454E4E53;
        16'h14E8 : rd_rsp_data <= 32'h804A5246;
        16'h14EC : rd_rsp_data <= 32'h80808080;
        16'h14F0 : rd_rsp_data <= 32'h80808080;
        16'h14F4 : rd_rsp_data <= 32'h014AA355;
        16'h14F8 : rd_rsp_data <= 32'h01020FFF;
        16'h14FC : rd_rsp_data <= 32'h01020FFF;
        16'h1500 : rd_rsp_data <= 32'h01020FFF;
        16'h1508 : rd_rsp_data <= 32'h001C937D;
        16'h150C : rd_rsp_data <= 32'h00FFFFFF;
        16'h1510 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1514 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1528 : rd_rsp_data <= 32'h03800000;
        16'h152C : rd_rsp_data <= 32'h070D19EE;
        16'h153C : rd_rsp_data <= 32'h023000E5;
        16'h1540 : rd_rsp_data <= 32'h0006087E;
        16'h1548 : rd_rsp_data <= 32'h80100010;
        16'h154C : rd_rsp_data <= 32'h99999999;
        16'h1550 : rd_rsp_data <= 32'h210841F0;
        16'h1554 : rd_rsp_data <= 32'h210842D0;
        16'h1558 : rd_rsp_data <= 32'h21084250;
        16'h155C : rd_rsp_data <= 32'h21084270;
        16'h1560 : rd_rsp_data <= 32'h21084210;
        16'h1564 : rd_rsp_data <= 32'h21084290;
        16'h1568 : rd_rsp_data <= 32'h21084230;
        16'h156C : rd_rsp_data <= 32'h210841F0;
        16'h1570 : rd_rsp_data <= 32'h21084210;
        16'h1574 : rd_rsp_data <= 32'h21084210;
        16'h1578 : rd_rsp_data <= 32'h00084210;
        16'h157C : rd_rsp_data <= 32'h00077054;
        16'h1580 : rd_rsp_data <= 32'h08400000;
        16'h1598 : rd_rsp_data <= 32'h808CF60A;
        16'h159C : rd_rsp_data <= 32'h00000016;
        16'h15A0 : rd_rsp_data <= 32'h00019400;
        16'h15AC : rd_rsp_data <= 32'h03260244;
        16'h15B0 : rd_rsp_data <= 32'h12481000;
        16'h15B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h15B8 : rd_rsp_data <= 32'h05800035;
        16'h15BC : rd_rsp_data <= 32'h0154C222;
        16'h15C4 : rd_rsp_data <= 32'h000003F6;
        16'h15C8 : rd_rsp_data <= 32'h78000000;
        16'h15D8 : rd_rsp_data <= 32'h07400000;
        16'h15DC : rd_rsp_data <= 32'h02180080;
        16'h15E0 : rd_rsp_data <= 32'h00162000;
        16'h15E8 : rd_rsp_data <= 32'h40000000;
        16'h1600 : rd_rsp_data <= 32'h00360C08;
        16'h1604 : rd_rsp_data <= 32'h00240808;
        16'h1608 : rd_rsp_data <= 32'h00101008;
        16'h160C : rd_rsp_data <= 32'h0035080C;
        16'h1610 : rd_rsp_data <= 32'h00140C0C;
        16'h1614 : rd_rsp_data <= 32'h00251410;
        16'h1618 : rd_rsp_data <= 32'h00200808;
        16'h161C : rd_rsp_data <= 32'h00240C0C;
        16'h1680 : rd_rsp_data <= 32'h10C68000;
        16'h1684 : rd_rsp_data <= 32'hF0783801;
        16'h1688 : rd_rsp_data <= 32'hFC212480;
        16'h168C : rd_rsp_data <= 32'h005D8001;
        16'h1690 : rd_rsp_data <= 32'h4F9E1000;
        16'h1694 : rd_rsp_data <= 32'h00063C21;
        16'h1698 : rd_rsp_data <= 32'h4DC00000;
        16'h169C : rd_rsp_data <= 32'h0A025B81;
        16'h16A0 : rd_rsp_data <= 32'h9FF057FE;
        16'h16A4 : rd_rsp_data <= 32'h7C210F7F;
        16'h16A8 : rd_rsp_data <= 32'h98C011DF;
        16'h16AC : rd_rsp_data <= 32'hA8000000;
        16'h16B0 : rd_rsp_data <= 32'h045E4904;
        16'h16B4 : rd_rsp_data <= 32'h061C003B;
        16'h16B8 : rd_rsp_data <= 32'h8820E21F;
        16'h16BC : rd_rsp_data <= 32'h58155D63;
        16'h16C8 : rd_rsp_data <= 32'h30000000;
        16'h16D4 : rd_rsp_data <= 32'h01041041;
        16'h16D8 : rd_rsp_data <= 32'h08208080;
        16'h16DC : rd_rsp_data <= 32'h1E560820;
        16'h16E0 : rd_rsp_data <= 32'h8062678C;
        16'h16E4 : rd_rsp_data <= 32'h5C6A645B;
        16'h16E8 : rd_rsp_data <= 32'h805E6751;
        16'h16EC : rd_rsp_data <= 32'h80808080;
        16'h16F0 : rd_rsp_data <= 32'h80808080;
        16'h16F4 : rd_rsp_data <= 32'h014292AB;
        16'h16F8 : rd_rsp_data <= 32'h01020FFF;
        16'h16FC : rd_rsp_data <= 32'h01020FFF;
        16'h1700 : rd_rsp_data <= 32'h01020FFF;
        16'h1708 : rd_rsp_data <= 32'h001C9379;
        16'h170C : rd_rsp_data <= 32'h00FFFFFF;
        16'h1710 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1714 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1720 : rd_rsp_data <= 32'h00003000;
        16'h1728 : rd_rsp_data <= 32'h03800000;
        16'h172C : rd_rsp_data <= 32'h074C1D7C;
        16'h173C : rd_rsp_data <= 32'h024604DC;
        16'h1740 : rd_rsp_data <= 32'h0006087E;
        16'h1748 : rd_rsp_data <= 32'h80100010;
        16'h174C : rd_rsp_data <= 32'h99999999;
        16'h1750 : rd_rsp_data <= 32'h21084230;
        16'h1754 : rd_rsp_data <= 32'h210841D0;
        16'h1758 : rd_rsp_data <= 32'h21084330;
        16'h175C : rd_rsp_data <= 32'h21084210;
        16'h1760 : rd_rsp_data <= 32'h210841F0;
        16'h1764 : rd_rsp_data <= 32'h21084250;
        16'h1768 : rd_rsp_data <= 32'h21084250;
        16'h176C : rd_rsp_data <= 32'h21084230;
        16'h1770 : rd_rsp_data <= 32'h21084210;
        16'h1774 : rd_rsp_data <= 32'h21084210;
        16'h1778 : rd_rsp_data <= 32'h00084210;
        16'h177C : rd_rsp_data <= 32'h00077054;
        16'h1780 : rd_rsp_data <= 32'h08400000;
        16'h1798 : rd_rsp_data <= 32'h808CF60A;
        16'h179C : rd_rsp_data <= 32'h00000016;
        16'h17A0 : rd_rsp_data <= 32'h00019400;
        16'h17AC : rd_rsp_data <= 32'h03260244;
        16'h17B0 : rd_rsp_data <= 32'h12481000;
        16'h17B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h17B8 : rd_rsp_data <= 32'h05800035;
        16'h17BC : rd_rsp_data <= 32'h0154C222;
        16'h17C4 : rd_rsp_data <= 32'h000007EC;
        16'h17C8 : rd_rsp_data <= 32'h7FF80000;
        16'h17D8 : rd_rsp_data <= 32'h07400000;
        16'h17DC : rd_rsp_data <= 32'h02180080;
        16'h17E0 : rd_rsp_data <= 32'h00162000;
        16'h17E8 : rd_rsp_data <= 32'h40000000;
        16'h1800 : rd_rsp_data <= 32'h00290C0C;
        16'h1804 : rd_rsp_data <= 32'h002D1D18;
        16'h1808 : rd_rsp_data <= 32'h00420C08;
        16'h180C : rd_rsp_data <= 32'h00141410;
        16'h1810 : rd_rsp_data <= 32'h002D1008;
        16'h1814 : rd_rsp_data <= 32'h00102519;
        16'h1818 : rd_rsp_data <= 32'h00211918;
        16'h181C : rd_rsp_data <= 32'h00292919;
        16'h1880 : rd_rsp_data <= 32'h10C68000;
        16'h1884 : rd_rsp_data <= 32'hF0F87843;
        16'h1888 : rd_rsp_data <= 32'hFC212480;
        16'h188C : rd_rsp_data <= 32'h005D0001;
        16'h1890 : rd_rsp_data <= 32'h4F9C1000;
        16'h1894 : rd_rsp_data <= 32'h00063C21;
        16'h1898 : rd_rsp_data <= 32'h4DE00000;
        16'h189C : rd_rsp_data <= 32'h0A025B81;
        16'h18A0 : rd_rsp_data <= 32'h9FF057FE;
        16'h18A4 : rd_rsp_data <= 32'hAC210FFB;
        16'h18A8 : rd_rsp_data <= 32'h98C011DF;
        16'h18AC : rd_rsp_data <= 32'hA8000000;
        16'h18B0 : rd_rsp_data <= 32'h045E4904;
        16'h18B4 : rd_rsp_data <= 32'h061C003B;
        16'h18B8 : rd_rsp_data <= 32'h8820EE1F;
        16'h18BC : rd_rsp_data <= 32'h58155D63;
        16'h18C8 : rd_rsp_data <= 32'h30000000;
        16'h18D4 : rd_rsp_data <= 32'h01041041;
        16'h18D8 : rd_rsp_data <= 32'h08208080;
        16'h18DC : rd_rsp_data <= 32'h1E560820;
        16'h18E0 : rd_rsp_data <= 32'h806B5E92;
        16'h18E4 : rd_rsp_data <= 32'h746C6C5E;
        16'h18E8 : rd_rsp_data <= 32'h805A745F;
        16'h18EC : rd_rsp_data <= 32'h80808080;
        16'h18F0 : rd_rsp_data <= 32'h80808080;
        16'h18F4 : rd_rsp_data <= 32'h016303A5;
        16'h18F8 : rd_rsp_data <= 32'h01020FFF;
        16'h18FC : rd_rsp_data <= 32'h01020FFF;
        16'h1900 : rd_rsp_data <= 32'h01020FFF;
        16'h1908 : rd_rsp_data <= 32'h002053A3;
        16'h190C : rd_rsp_data <= 32'h00FFFFFF;
        16'h1910 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1914 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1920 : rd_rsp_data <= 32'h00003000;
        16'h1928 : rd_rsp_data <= 32'h03800000;
        16'h192C : rd_rsp_data <= 32'h0640BFA5;
        16'h193C : rd_rsp_data <= 32'h023404E3;
        16'h1940 : rd_rsp_data <= 32'h0006087E;
        16'h1948 : rd_rsp_data <= 32'h80100010;
        16'h194C : rd_rsp_data <= 32'h99999999;
        16'h1950 : rd_rsp_data <= 32'h210841F0;
        16'h1954 : rd_rsp_data <= 32'h21084250;
        16'h1958 : rd_rsp_data <= 32'h21084290;
        16'h195C : rd_rsp_data <= 32'h21084290;
        16'h1960 : rd_rsp_data <= 32'h21084210;
        16'h1964 : rd_rsp_data <= 32'h21084230;
        16'h1968 : rd_rsp_data <= 32'h21084210;
        16'h196C : rd_rsp_data <= 32'h21084230;
        16'h1970 : rd_rsp_data <= 32'h21084210;
        16'h1974 : rd_rsp_data <= 32'h21084210;
        16'h1978 : rd_rsp_data <= 32'h00084210;
        16'h197C : rd_rsp_data <= 32'h00077054;
        16'h1980 : rd_rsp_data <= 32'h08400000;
        16'h1998 : rd_rsp_data <= 32'h808CF60A;
        16'h199C : rd_rsp_data <= 32'h00000010;
        16'h19A0 : rd_rsp_data <= 32'h00019400;
        16'h19AC : rd_rsp_data <= 32'h03260244;
        16'h19B0 : rd_rsp_data <= 32'h12481000;
        16'h19B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h19B8 : rd_rsp_data <= 32'h05800035;
        16'h19BC : rd_rsp_data <= 32'h0154C222;
        16'h19C4 : rd_rsp_data <= 32'h000006BE;
        16'h19C8 : rd_rsp_data <= 32'h78000000;
        16'h19D8 : rd_rsp_data <= 32'h07400000;
        16'h19DC : rd_rsp_data <= 32'h02180080;
        16'h19E0 : rd_rsp_data <= 32'h00102000;
        16'h19E8 : rd_rsp_data <= 32'h40000000;
        16'h1A00 : rd_rsp_data <= 32'h0025140C;
        16'h1A04 : rd_rsp_data <= 32'h002D1008;
        16'h1A08 : rd_rsp_data <= 32'h003A1410;
        16'h1A0C : rd_rsp_data <= 32'h0014140C;
        16'h1A10 : rd_rsp_data <= 32'h00081D14;
        16'h1A14 : rd_rsp_data <= 32'h00291008;
        16'h1A18 : rd_rsp_data <= 32'h00201C15;
        16'h1A1C : rd_rsp_data <= 32'h00251008;
        16'h1A80 : rd_rsp_data <= 32'h10C68000;
        16'h1A84 : rd_rsp_data <= 32'hF0F87843;
        16'h1A88 : rd_rsp_data <= 32'hFC212480;
        16'h1A8C : rd_rsp_data <= 32'h005E4001;
        16'h1A90 : rd_rsp_data <= 32'h4F1E1000;
        16'h1A94 : rd_rsp_data <= 32'h00063C21;
        16'h1A98 : rd_rsp_data <= 32'h55E00000;
        16'h1A9C : rd_rsp_data <= 32'h0A025B81;
        16'h1AA0 : rd_rsp_data <= 32'h9FF056BE;
        16'h1AA4 : rd_rsp_data <= 32'h7C210FF9;
        16'h1AA8 : rd_rsp_data <= 32'h98C011DF;
        16'h1AAC : rd_rsp_data <= 32'hA8000000;
        16'h1AB0 : rd_rsp_data <= 32'h045E4904;
        16'h1AB4 : rd_rsp_data <= 32'h061C003B;
        16'h1AB8 : rd_rsp_data <= 32'h8820E21F;
        16'h1ABC : rd_rsp_data <= 32'h58155D63;
        16'h1AC8 : rd_rsp_data <= 32'h30000000;
        16'h1AD4 : rd_rsp_data <= 32'h01041041;
        16'h1AD8 : rd_rsp_data <= 32'h08208080;
        16'h1ADC : rd_rsp_data <= 32'h1E560820;
        16'h1AE0 : rd_rsp_data <= 32'h805C50A3;
        16'h1AE4 : rd_rsp_data <= 32'h59575C50;
        16'h1AE8 : rd_rsp_data <= 32'h804E524A;
        16'h1AEC : rd_rsp_data <= 32'h80808080;
        16'h1AF0 : rd_rsp_data <= 32'h80808080;
        16'h1AF4 : rd_rsp_data <= 32'h016B130B;
        16'h1AF8 : rd_rsp_data <= 32'h01020FFF;
        16'h1AFC : rd_rsp_data <= 32'h01020FFF;
        16'h1B00 : rd_rsp_data <= 32'h01020FFF;
        16'h1B08 : rd_rsp_data <= 32'h0021D3BD;
        16'h1B0C : rd_rsp_data <= 32'h00FFFFFF;
        16'h1B10 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1B14 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1B20 : rd_rsp_data <= 32'h00003000;
        16'h1B28 : rd_rsp_data <= 32'h03800000;
        16'h1B2C : rd_rsp_data <= 32'h0640BBBC;
        16'h1B3C : rd_rsp_data <= 32'h023A00E1;
        16'h1B40 : rd_rsp_data <= 32'h0006087E;
        16'h1B48 : rd_rsp_data <= 32'h80100010;
        16'h1B4C : rd_rsp_data <= 32'h99999999;
        16'h1B50 : rd_rsp_data <= 32'h21084230;
        16'h1B54 : rd_rsp_data <= 32'h21084210;
        16'h1B58 : rd_rsp_data <= 32'h210841F0;
        16'h1B5C : rd_rsp_data <= 32'h21084230;
        16'h1B60 : rd_rsp_data <= 32'h21084290;
        16'h1B64 : rd_rsp_data <= 32'h210841D0;
        16'h1B68 : rd_rsp_data <= 32'h21084210;
        16'h1B6C : rd_rsp_data <= 32'h21084210;
        16'h1B70 : rd_rsp_data <= 32'h21084210;
        16'h1B74 : rd_rsp_data <= 32'h21084210;
        16'h1B78 : rd_rsp_data <= 32'h00084210;
        16'h1B7C : rd_rsp_data <= 32'h00077054;
        16'h1B80 : rd_rsp_data <= 32'h08400000;
        16'h1B98 : rd_rsp_data <= 32'h808CF60A;
        16'h1B9C : rd_rsp_data <= 32'h00000018;
        16'h1BA0 : rd_rsp_data <= 32'h00019400;
        16'h1BAC : rd_rsp_data <= 32'h03260244;
        16'h1BB0 : rd_rsp_data <= 32'h12481000;
        16'h1BB4 : rd_rsp_data <= 32'h2D495C3E;
        16'h1BB8 : rd_rsp_data <= 32'h05800035;
        16'h1BBC : rd_rsp_data <= 32'h0154C222;
        16'h1BC4 : rd_rsp_data <= 32'h000005DE;
        16'h1BC8 : rd_rsp_data <= 32'h78000000;
        16'h1BD8 : rd_rsp_data <= 32'h07400000;
        16'h1BDC : rd_rsp_data <= 32'h02180080;
        16'h1BE0 : rd_rsp_data <= 32'h00182000;
        16'h1BE8 : rd_rsp_data <= 32'h40000000;
        16'h1C00 : rd_rsp_data <= 32'h00241D21;
        16'h1C04 : rd_rsp_data <= 32'h0031100C;
        16'h1C08 : rd_rsp_data <= 32'h00181419;
        16'h1C0C : rd_rsp_data <= 32'h002C100C;
        16'h1C10 : rd_rsp_data <= 32'h00281410;
        16'h1C14 : rd_rsp_data <= 32'h0042100C;
        16'h1C18 : rd_rsp_data <= 32'h0028100C;
        16'h1C1C : rd_rsp_data <= 32'h00420C08;
        16'h1C80 : rd_rsp_data <= 32'h10C68000;
        16'h1C84 : rd_rsp_data <= 32'hF0F87843;
        16'h1C88 : rd_rsp_data <= 32'hFC212480;
        16'h1C8C : rd_rsp_data <= 32'h00590001;
        16'h1C90 : rd_rsp_data <= 32'h4F1E1000;
        16'h1C94 : rd_rsp_data <= 32'h00063C21;
        16'h1C98 : rd_rsp_data <= 32'h5DE00000;
        16'h1C9C : rd_rsp_data <= 32'h0A025B81;
        16'h1CA0 : rd_rsp_data <= 32'h9FF056BE;
        16'h1CA4 : rd_rsp_data <= 32'h9C210F7C;
        16'h1CA8 : rd_rsp_data <= 32'h98C011DF;
        16'h1CAC : rd_rsp_data <= 32'hA8000000;
        16'h1CB0 : rd_rsp_data <= 32'h045E4904;
        16'h1CB4 : rd_rsp_data <= 32'h061C003B;
        16'h1CB8 : rd_rsp_data <= 32'h8820F21F;
        16'h1CBC : rd_rsp_data <= 32'h58155D63;
        16'h1CC8 : rd_rsp_data <= 32'h30000000;
        16'h1CD4 : rd_rsp_data <= 32'h01041041;
        16'h1CD8 : rd_rsp_data <= 32'h08208080;
        16'h1CDC : rd_rsp_data <= 32'h1E560820;
        16'h1CE0 : rd_rsp_data <= 32'h80666888;
        16'h1CE4 : rd_rsp_data <= 32'h685E5A70;
        16'h1CE8 : rd_rsp_data <= 32'h805C615D;
        16'h1CEC : rd_rsp_data <= 32'h80808080;
        16'h1CF0 : rd_rsp_data <= 32'h80808080;
        16'h1CF4 : rd_rsp_data <= 32'h018323B5;
        16'h1CF8 : rd_rsp_data <= 32'h01020FFF;
        16'h1CFC : rd_rsp_data <= 32'h01020FFF;
        16'h1D00 : rd_rsp_data <= 32'h01020FFF;
        16'h1D08 : rd_rsp_data <= 32'h001FD3A1;
        16'h1D0C : rd_rsp_data <= 32'h00FFFFFF;
        16'h1D10 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1D14 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1D28 : rd_rsp_data <= 32'h03800000;
        16'h1D2C : rd_rsp_data <= 32'h0740BFA5;
        16'h1D3C : rd_rsp_data <= 32'h023404E3;
        16'h1D40 : rd_rsp_data <= 32'h0006087E;
        16'h1D48 : rd_rsp_data <= 32'h80100010;
        16'h1D4C : rd_rsp_data <= 32'h99999999;
        16'h1D50 : rd_rsp_data <= 32'h210842B0;
        16'h1D54 : rd_rsp_data <= 32'h21084270;
        16'h1D58 : rd_rsp_data <= 32'h210841F0;
        16'h1D5C : rd_rsp_data <= 32'h210842B0;
        16'h1D60 : rd_rsp_data <= 32'h21084250;
        16'h1D64 : rd_rsp_data <= 32'h210842B0;
        16'h1D68 : rd_rsp_data <= 32'h210842B0;
        16'h1D6C : rd_rsp_data <= 32'h21084290;
        16'h1D70 : rd_rsp_data <= 32'h21084210;
        16'h1D74 : rd_rsp_data <= 32'h21084210;
        16'h1D78 : rd_rsp_data <= 32'h00084210;
        16'h1D7C : rd_rsp_data <= 32'h00077054;
        16'h1D80 : rd_rsp_data <= 32'h08400000;
        16'h1D98 : rd_rsp_data <= 32'h808CF60A;
        16'h1D9C : rd_rsp_data <= 32'h00000016;
        16'h1DA0 : rd_rsp_data <= 32'h00019400;
        16'h1DAC : rd_rsp_data <= 32'h03260244;
        16'h1DB0 : rd_rsp_data <= 32'h12481000;
        16'h1DB4 : rd_rsp_data <= 32'h2D495C3E;
        16'h1DB8 : rd_rsp_data <= 32'h05800035;
        16'h1DBC : rd_rsp_data <= 32'h0154C222;
        16'h1DC4 : rd_rsp_data <= 32'h000000BC;
        16'h1DC8 : rd_rsp_data <= 32'h78000000;
        16'h1DD8 : rd_rsp_data <= 32'h07400000;
        16'h1DDC : rd_rsp_data <= 32'h02180080;
        16'h1DE0 : rd_rsp_data <= 32'h00162000;
        16'h1DE8 : rd_rsp_data <= 32'h40000000;
        16'h1E00 : rd_rsp_data <= 32'h00252A20;
        16'h1E04 : rd_rsp_data <= 32'h00183229;
        16'h1E08 : rd_rsp_data <= 32'h000C2514;
        16'h1E0C : rd_rsp_data <= 32'h0010251D;
        16'h1E10 : rd_rsp_data <= 32'h00102118;
        16'h1E14 : rd_rsp_data <= 32'h00202114;
        16'h1E18 : rd_rsp_data <= 32'h002D140C;
        16'h1E1C : rd_rsp_data <= 32'h00322118;
        16'h1E80 : rd_rsp_data <= 32'h10C68000;
        16'h1E84 : rd_rsp_data <= 32'hF0F87843;
        16'h1E88 : rd_rsp_data <= 32'hFC212480;
        16'h1E8C : rd_rsp_data <= 32'h0059C001;
        16'h1E90 : rd_rsp_data <= 32'h4E1E1000;
        16'h1E94 : rd_rsp_data <= 32'h00063C21;
        16'h1E98 : rd_rsp_data <= 32'h46800000;
        16'h1E9C : rd_rsp_data <= 32'h0A025B81;
        16'h1EA0 : rd_rsp_data <= 32'h9FF057BE;
        16'h1EA4 : rd_rsp_data <= 32'h14210F9F;
        16'h1EA8 : rd_rsp_data <= 32'h98C011DF;
        16'h1EAC : rd_rsp_data <= 32'hA8000000;
        16'h1EB0 : rd_rsp_data <= 32'h045E4904;
        16'h1EB4 : rd_rsp_data <= 32'h061C003B;
        16'h1EB8 : rd_rsp_data <= 32'h8820EE1F;
        16'h1EBC : rd_rsp_data <= 32'h58155D63;
        16'h1EC8 : rd_rsp_data <= 32'h30000000;
        16'h1ED4 : rd_rsp_data <= 32'h01041041;
        16'h1ED8 : rd_rsp_data <= 32'h08208080;
        16'h1EDC : rd_rsp_data <= 32'h1E560820;
        16'h1EE0 : rd_rsp_data <= 32'h80584E93;
        16'h1EE4 : rd_rsp_data <= 32'h52605562;
        16'h1EE8 : rd_rsp_data <= 32'h805B5C4A;
        16'h1EEC : rd_rsp_data <= 32'h80808080;
        16'h1EF0 : rd_rsp_data <= 32'h80808080;
        16'h1EF4 : rd_rsp_data <= 32'h0142E323;
        16'h1EF8 : rd_rsp_data <= 32'h01020FFF;
        16'h1EFC : rd_rsp_data <= 32'h01020FFF;
        16'h1F00 : rd_rsp_data <= 32'h01020FFF;
        16'h1F08 : rd_rsp_data <= 32'h002093B3;
        16'h1F0C : rd_rsp_data <= 32'h00FFFFFF;
        16'h1F10 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1F14 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1F20 : rd_rsp_data <= 32'h0001D000;
        16'h1F28 : rd_rsp_data <= 32'h03800000;
        16'h1F2C : rd_rsp_data <= 32'h0740BBBC;
        16'h1F3C : rd_rsp_data <= 32'h023A00E1;
        16'h1F40 : rd_rsp_data <= 32'h0006087E;
        16'h1F48 : rd_rsp_data <= 32'h80100010;
        16'h1F4C : rd_rsp_data <= 32'h99999999;
        16'h1F50 : rd_rsp_data <= 32'h21084190;
        16'h1F54 : rd_rsp_data <= 32'h21084190;
        16'h1F58 : rd_rsp_data <= 32'h210841F0;
        16'h1F5C : rd_rsp_data <= 32'h21084230;
        16'h1F60 : rd_rsp_data <= 32'h21084290;
        16'h1F64 : rd_rsp_data <= 32'h210842B0;
        16'h1F68 : rd_rsp_data <= 32'h210841D0;
        16'h1F6C : rd_rsp_data <= 32'h21084210;
        16'h1F70 : rd_rsp_data <= 32'h21084210;
        16'h1F74 : rd_rsp_data <= 32'h21084210;
        16'h1F78 : rd_rsp_data <= 32'h00084210;
        16'h1F7C : rd_rsp_data <= 32'h00077054;
        16'h1F80 : rd_rsp_data <= 32'h08400000;
        16'h1F98 : rd_rsp_data <= 32'h808CF60A;
        16'h1F9C : rd_rsp_data <= 32'h00000018;
        16'h1FA0 : rd_rsp_data <= 32'h00019400;
        16'h1FAC : rd_rsp_data <= 32'h03260244;
        16'h1FB0 : rd_rsp_data <= 32'h12481000;
        16'h1FB4 : rd_rsp_data <= 32'h2D495C3E;
        16'h1FB8 : rd_rsp_data <= 32'h05800035;
        16'h1FBC : rd_rsp_data <= 32'h0154C222;
        16'h1FC4 : rd_rsp_data <= 32'h0000014E;
        16'h1FC8 : rd_rsp_data <= 32'h78000000;
        16'h1FD8 : rd_rsp_data <= 32'h07400000;
        16'h1FDC : rd_rsp_data <= 32'h02180080;
        16'h1FE0 : rd_rsp_data <= 32'h00182000;
        16'h1FE8 : rd_rsp_data <= 32'h40000000;
        16'h2080 : rd_rsp_data <= 32'h010600A0;
        16'h2088 : rd_rsp_data <= 32'hBC012400;
        16'h208C : rd_rsp_data <= 32'h00400000;
        16'h2090 : rd_rsp_data <= 32'h0C4A1800;
        16'h2094 : rd_rsp_data <= 32'h00043C42;
        16'h2098 : rd_rsp_data <= 32'h0C200000;
        16'h209C : rd_rsp_data <= 32'h00038381;
        16'h20A0 : rd_rsp_data <= 32'h187037FE;
        16'h20A4 : rd_rsp_data <= 32'h84210FFF;
        16'h20A8 : rd_rsp_data <= 32'hC00011C3;
        16'h20B0 : rd_rsp_data <= 32'h00002904;
        16'h20B4 : rd_rsp_data <= 32'h061D0238;
        16'h20B8 : rd_rsp_data <= 32'h0820221A;
        16'h20BC : rd_rsp_data <= 32'h0813A0A4;
        16'h20C8 : rd_rsp_data <= 32'h38000000;
        16'h20D4 : rd_rsp_data <= 32'h01041040;
        16'h20D8 : rd_rsp_data <= 32'h08201010;
        16'h20DC : rd_rsp_data <= 32'h203A0820;
        16'h20E0 : rd_rsp_data <= 32'h80808080;
        16'h20E4 : rd_rsp_data <= 32'h80808080;
        16'h20E8 : rd_rsp_data <= 32'h80808080;
        16'h20EC : rd_rsp_data <= 32'h80808080;
        16'h20F0 : rd_rsp_data <= 32'h80808080;
        16'h20F4 : rd_rsp_data <= 32'h01020FFF;
        16'h20F8 : rd_rsp_data <= 32'h01020FFF;
        16'h20FC : rd_rsp_data <= 32'h01020FFF;
        16'h2100 : rd_rsp_data <= 32'h01020FFF;
        16'h2108 : rd_rsp_data <= 32'h00FFFFFF;
        16'h210C : rd_rsp_data <= 32'h00FFFFFF;
        16'h2110 : rd_rsp_data <= 32'h00FFFFFF;
        16'h2114 : rd_rsp_data <= 32'h00FFFFFF;
        16'h212C : rd_rsp_data <= 32'h00FAC688;
        16'h2148 : rd_rsp_data <= 32'h80100000;
        16'h214C : rd_rsp_data <= 32'h88888888;
        16'h2150 : rd_rsp_data <= 32'h21084210;
        16'h2154 : rd_rsp_data <= 32'h21084210;
        16'h2158 : rd_rsp_data <= 32'h21084210;
        16'h215C : rd_rsp_data <= 32'h21084210;
        16'h2160 : rd_rsp_data <= 32'h21084210;
        16'h2164 : rd_rsp_data <= 32'h21084210;
        16'h2168 : rd_rsp_data <= 32'h21084210;
        16'h216C : rd_rsp_data <= 32'h21084210;
        16'h2170 : rd_rsp_data <= 32'h21084210;
        16'h2174 : rd_rsp_data <= 32'h21084210;
        16'h2178 : rd_rsp_data <= 32'h00084210;
        16'h217C : rd_rsp_data <= 32'h00024254;
        16'h2180 : rd_rsp_data <= 32'h08400000;
        16'h219C : rd_rsp_data <= 32'h00000400;
        16'h21AC : rd_rsp_data <= 32'h03260244;
        16'h21B0 : rd_rsp_data <= 32'h12481000;
        16'h21B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h21B8 : rd_rsp_data <= 32'h05800035;
        16'h21BC : rd_rsp_data <= 32'h0154C222;
        16'h21C4 : rd_rsp_data <= 32'h000002DE;
        16'h21C8 : rd_rsp_data <= 32'h78000000;
        16'h21D8 : rd_rsp_data <= 32'h02000000;
        16'h21DC : rd_rsp_data <= 32'h02180080;
        16'h21E0 : rd_rsp_data <= 32'h00002000;
        16'h21E8 : rd_rsp_data <= 32'h40000000;
        16'h2280 : rd_rsp_data <= 32'h010600A0;
        16'h2288 : rd_rsp_data <= 32'hBC012400;
        16'h228C : rd_rsp_data <= 32'h00400000;
        16'h2290 : rd_rsp_data <= 32'h0C4A1800;
        16'h2294 : rd_rsp_data <= 32'h00043C42;
        16'h2298 : rd_rsp_data <= 32'h0C200000;
        16'h229C : rd_rsp_data <= 32'h00038381;
        16'h22A0 : rd_rsp_data <= 32'h187037FE;
        16'h22A4 : rd_rsp_data <= 32'h84210FFF;
        16'h22A8 : rd_rsp_data <= 32'hC00011C3;
        16'h22B0 : rd_rsp_data <= 32'h00002904;
        16'h22B4 : rd_rsp_data <= 32'h061D0238;
        16'h22B8 : rd_rsp_data <= 32'h0820221A;
        16'h22BC : rd_rsp_data <= 32'h0813A0A4;
        16'h22C8 : rd_rsp_data <= 32'h38000000;
        16'h22D4 : rd_rsp_data <= 32'h01041040;
        16'h22D8 : rd_rsp_data <= 32'h08201010;
        16'h22DC : rd_rsp_data <= 32'h203A0820;
        16'h22E0 : rd_rsp_data <= 32'h80808080;
        16'h22E4 : rd_rsp_data <= 32'h80808080;
        16'h22E8 : rd_rsp_data <= 32'h80808080;
        16'h22EC : rd_rsp_data <= 32'h80808080;
        16'h22F0 : rd_rsp_data <= 32'h80808080;
        16'h22F4 : rd_rsp_data <= 32'h01020FFF;
        16'h22F8 : rd_rsp_data <= 32'h01020FFF;
        16'h22FC : rd_rsp_data <= 32'h01020FFF;
        16'h2300 : rd_rsp_data <= 32'h01020FFF;
        16'h2308 : rd_rsp_data <= 32'h00FFFFFF;
        16'h230C : rd_rsp_data <= 32'h00FFFFFF;
        16'h2310 : rd_rsp_data <= 32'h00FFFFFF;
        16'h2314 : rd_rsp_data <= 32'h00FFFFFF;
        16'h232C : rd_rsp_data <= 32'h00FAC688;
        16'h2348 : rd_rsp_data <= 32'h80100000;
        16'h234C : rd_rsp_data <= 32'h88888888;
        16'h2350 : rd_rsp_data <= 32'h21084210;
        16'h2354 : rd_rsp_data <= 32'h21084210;
        16'h2358 : rd_rsp_data <= 32'h21084210;
        16'h235C : rd_rsp_data <= 32'h21084210;
        16'h2360 : rd_rsp_data <= 32'h21084210;
        16'h2364 : rd_rsp_data <= 32'h21084210;
        16'h2368 : rd_rsp_data <= 32'h21084210;
        16'h236C : rd_rsp_data <= 32'h21084210;
        16'h2370 : rd_rsp_data <= 32'h21084210;
        16'h2374 : rd_rsp_data <= 32'h21084210;
        16'h2378 : rd_rsp_data <= 32'h00084210;
        16'h237C : rd_rsp_data <= 32'h00024254;
        16'h2380 : rd_rsp_data <= 32'h08400000;
        16'h239C : rd_rsp_data <= 32'h00000400;
        16'h23AC : rd_rsp_data <= 32'h03260244;
        16'h23B0 : rd_rsp_data <= 32'h12481000;
        16'h23B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h23B8 : rd_rsp_data <= 32'h05800035;
        16'h23BC : rd_rsp_data <= 32'h0154C222;
        16'h23C4 : rd_rsp_data <= 32'h000003D6;
        16'h23C8 : rd_rsp_data <= 32'h78000000;
        16'h23D8 : rd_rsp_data <= 32'h02000000;
        16'h23DC : rd_rsp_data <= 32'h02180080;
        16'h23E0 : rd_rsp_data <= 32'h00002000;
        16'h23E8 : rd_rsp_data <= 32'h40000000;
        16'h2480 : rd_rsp_data <= 32'h010600A0;
        16'h2488 : rd_rsp_data <= 32'hBC012400;
        16'h248C : rd_rsp_data <= 32'h00400000;
        16'h2490 : rd_rsp_data <= 32'h0C4A1800;
        16'h2494 : rd_rsp_data <= 32'h00043C42;
        16'h2498 : rd_rsp_data <= 32'h0C200000;
        16'h249C : rd_rsp_data <= 32'h00038381;
        16'h24A0 : rd_rsp_data <= 32'h187037FE;
        16'h24A4 : rd_rsp_data <= 32'h84210FFF;
        16'h24A8 : rd_rsp_data <= 32'hC00011C3;
        16'h24B0 : rd_rsp_data <= 32'h00002904;
        16'h24B4 : rd_rsp_data <= 32'h061D0238;
        16'h24B8 : rd_rsp_data <= 32'h0820221A;
        16'h24BC : rd_rsp_data <= 32'h0813A0A4;
        16'h24C8 : rd_rsp_data <= 32'h38000000;
        16'h24D4 : rd_rsp_data <= 32'h01041040;
        16'h24D8 : rd_rsp_data <= 32'h08201010;
        16'h24DC : rd_rsp_data <= 32'h203A0820;
        16'h24E0 : rd_rsp_data <= 32'h80808080;
        16'h24E4 : rd_rsp_data <= 32'h80808080;
        16'h24E8 : rd_rsp_data <= 32'h80808080;
        16'h24EC : rd_rsp_data <= 32'h80808080;
        16'h24F0 : rd_rsp_data <= 32'h80808080;
        16'h24F4 : rd_rsp_data <= 32'h01020FFF;
        16'h24F8 : rd_rsp_data <= 32'h01020FFF;
        16'h24FC : rd_rsp_data <= 32'h01020FFF;
        16'h2500 : rd_rsp_data <= 32'h01020FFF;
        16'h2508 : rd_rsp_data <= 32'h00FFFFFF;
        16'h250C : rd_rsp_data <= 32'h00FFFFFF;
        16'h2510 : rd_rsp_data <= 32'h00FFFFFF;
        16'h2514 : rd_rsp_data <= 32'h00FFFFFF;
        16'h252C : rd_rsp_data <= 32'h00FAC688;
        16'h2548 : rd_rsp_data <= 32'h80100000;
        16'h254C : rd_rsp_data <= 32'h88888888;
        16'h2550 : rd_rsp_data <= 32'h21084210;
        16'h2554 : rd_rsp_data <= 32'h21084210;
        16'h2558 : rd_rsp_data <= 32'h21084210;
        16'h255C : rd_rsp_data <= 32'h21084210;
        16'h2560 : rd_rsp_data <= 32'h21084210;
        16'h2564 : rd_rsp_data <= 32'h21084210;
        16'h2568 : rd_rsp_data <= 32'h21084210;
        16'h256C : rd_rsp_data <= 32'h21084210;
        16'h2570 : rd_rsp_data <= 32'h21084210;
        16'h2574 : rd_rsp_data <= 32'h21084210;
        16'h2578 : rd_rsp_data <= 32'h00084210;
        16'h257C : rd_rsp_data <= 32'h00024254;
        16'h2580 : rd_rsp_data <= 32'h08400000;
        16'h259C : rd_rsp_data <= 32'h00000400;
        16'h25AC : rd_rsp_data <= 32'h03260244;
        16'h25B0 : rd_rsp_data <= 32'h12481000;
        16'h25B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h25B8 : rd_rsp_data <= 32'h05800035;
        16'h25BC : rd_rsp_data <= 32'h0154C222;
        16'h25C4 : rd_rsp_data <= 32'h000007FE;
        16'h25C8 : rd_rsp_data <= 32'h78000000;
        16'h25D8 : rd_rsp_data <= 32'h02000000;
        16'h25DC : rd_rsp_data <= 32'h02180080;
        16'h25E0 : rd_rsp_data <= 32'h00002000;
        16'h25E8 : rd_rsp_data <= 32'h40000000;
        16'h2680 : rd_rsp_data <= 32'h010600A0;
        16'h2688 : rd_rsp_data <= 32'hBC012400;
        16'h268C : rd_rsp_data <= 32'h00400000;
        16'h2690 : rd_rsp_data <= 32'h0C4A1800;
        16'h2694 : rd_rsp_data <= 32'h00043C42;
        16'h2698 : rd_rsp_data <= 32'h0C200000;
        16'h269C : rd_rsp_data <= 32'h00038381;
        16'h26A0 : rd_rsp_data <= 32'h187037FE;
        16'h26A4 : rd_rsp_data <= 32'h84210FFF;
        16'h26A8 : rd_rsp_data <= 32'hC00011C3;
        16'h26B0 : rd_rsp_data <= 32'h00002904;
        16'h26B4 : rd_rsp_data <= 32'h061D0238;
        16'h26B8 : rd_rsp_data <= 32'h0820221A;
        16'h26BC : rd_rsp_data <= 32'h0813A0A4;
        16'h26C8 : rd_rsp_data <= 32'h38000000;
        16'h26D4 : rd_rsp_data <= 32'h01041040;
        16'h26D8 : rd_rsp_data <= 32'h08201010;
        16'h26DC : rd_rsp_data <= 32'h203A0820;
        16'h26E0 : rd_rsp_data <= 32'h80808080;
        16'h26E4 : rd_rsp_data <= 32'h80808080;
        16'h26E8 : rd_rsp_data <= 32'h80808080;
        16'h26EC : rd_rsp_data <= 32'h80808080;
        16'h26F0 : rd_rsp_data <= 32'h80808080;
        16'h26F4 : rd_rsp_data <= 32'h01020FFF;
        16'h26F8 : rd_rsp_data <= 32'h01020FFF;
        16'h26FC : rd_rsp_data <= 32'h01020FFF;
        16'h2700 : rd_rsp_data <= 32'h01020FFF;
        16'h2708 : rd_rsp_data <= 32'h00FFFFFF;
        16'h270C : rd_rsp_data <= 32'h00FFFFFF;
        16'h2710 : rd_rsp_data <= 32'h00FFFFFF;
        16'h2714 : rd_rsp_data <= 32'h00FFFFFF;
        16'h272C : rd_rsp_data <= 32'h00FAC688;
        16'h2748 : rd_rsp_data <= 32'h80100000;
        16'h274C : rd_rsp_data <= 32'h88888888;
        16'h2750 : rd_rsp_data <= 32'h21084210;
        16'h2754 : rd_rsp_data <= 32'h21084210;
        16'h2758 : rd_rsp_data <= 32'h21084210;
        16'h275C : rd_rsp_data <= 32'h21084210;
        16'h2760 : rd_rsp_data <= 32'h21084210;
        16'h2764 : rd_rsp_data <= 32'h21084210;
        16'h2768 : rd_rsp_data <= 32'h21084210;
        16'h276C : rd_rsp_data <= 32'h21084210;
        16'h2770 : rd_rsp_data <= 32'h21084210;
        16'h2774 : rd_rsp_data <= 32'h21084210;
        16'h2778 : rd_rsp_data <= 32'h00084210;
        16'h277C : rd_rsp_data <= 32'h00024254;
        16'h2780 : rd_rsp_data <= 32'h08400000;
        16'h279C : rd_rsp_data <= 32'h00000400;
        16'h27AC : rd_rsp_data <= 32'h03260244;
        16'h27B0 : rd_rsp_data <= 32'h12481000;
        16'h27B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h27B8 : rd_rsp_data <= 32'h05800035;
        16'h27BC : rd_rsp_data <= 32'h0154C222;
        16'h27C4 : rd_rsp_data <= 32'h000006E0;
        16'h27C8 : rd_rsp_data <= 32'h78000000;
        16'h27D8 : rd_rsp_data <= 32'h02000000;
        16'h27DC : rd_rsp_data <= 32'h02180080;
        16'h27E0 : rd_rsp_data <= 32'h00002000;
        16'h27E8 : rd_rsp_data <= 32'h40000000;
        16'h2800 : rd_rsp_data <= 32'h00001503;
        16'h2804 : rd_rsp_data <= 32'h00FF0F0F;
        16'h2808 : rd_rsp_data <= 32'h00082315;
        16'h2880 : rd_rsp_data <= 32'h00001503;
        16'h2884 : rd_rsp_data <= 32'h00FF0F0F;
        16'h2888 : rd_rsp_data <= 32'h00082315;
        16'h2900 : rd_rsp_data <= 32'h00000003;
        16'h2908 : rd_rsp_data <= 32'h0640E9A0;
        16'h2910 : rd_rsp_data <= 32'h3BF7EFBD;
        16'h2914 : rd_rsp_data <= 32'h0000003E;
        16'h2918 : rd_rsp_data <= 32'h00000001;
        16'h2980 : rd_rsp_data <= 32'h00000003;
        16'h2988 : rd_rsp_data <= 32'h0640E9A0;
        16'h2990 : rd_rsp_data <= 32'h3BF7FF3D;
        16'h2994 : rd_rsp_data <= 32'h0000003E;
        16'h2998 : rd_rsp_data <= 32'h00000001;
        16'h2A00 : rd_rsp_data <= 32'h00000003;
        16'h2A08 : rd_rsp_data <= 32'h0640E9A0;
        16'h2A10 : rd_rsp_data <= 32'h3DFBEF3F;
        16'h2A14 : rd_rsp_data <= 32'h0000003E;
        16'h2A18 : rd_rsp_data <= 32'h00000001;
        16'h2A80 : rd_rsp_data <= 32'h00000003;
        16'h2A88 : rd_rsp_data <= 32'h0640E9A0;
        16'h2A90 : rd_rsp_data <= 32'h3F03EF80;
        16'h2A98 : rd_rsp_data <= 32'h00000001;
        16'h2B00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2B9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2BFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h2C00 : rd_rsp_data <= 32'h0001860E;
        16'h2C04 : rd_rsp_data <= 32'h00015820;
        16'h2C0C : rd_rsp_data <= 32'h6C820008;
        16'h2C10 : rd_rsp_data <= 32'h00000402;
        16'h2C14 : rd_rsp_data <= 32'h3B000001;
        16'h2C18 : rd_rsp_data <= 32'hC1B20022;
        16'h2C1C : rd_rsp_data <= 32'h00410000;
        16'h2C20 : rd_rsp_data <= 32'h00000100;
        16'h2C24 : rd_rsp_data <= 32'h10003001;
        16'h2C28 : rd_rsp_data <= 32'h10100000;
        16'h2C2C : rd_rsp_data <= 32'h0010E2C0;
        16'h2C30 : rd_rsp_data <= 32'h1831BD44;
        16'h2C34 : rd_rsp_data <= 32'h0182B060;
        16'h2C38 : rd_rsp_data <= 32'hC0040534;
        16'h2C3C : rd_rsp_data <= 32'h602AD500;
        16'h2C40 : rd_rsp_data <= 32'hE0D50000;
        16'h2C48 : rd_rsp_data <= 32'h13004000;
        16'h2C4C : rd_rsp_data <= 32'h3C130E40;
        16'h2C50 : rd_rsp_data <= 32'h0145930E;
        16'h2C54 : rd_rsp_data <= 32'hFCD068AD;
        16'h2C58 : rd_rsp_data <= 32'h6C9B3062;
        16'h2C5C : rd_rsp_data <= 32'h00000001;
        16'h2C60 : rd_rsp_data <= 32'h1C104457;
        16'h2C64 : rd_rsp_data <= 32'h00006C82;
        16'h2C6C : rd_rsp_data <= 32'h04000000;
        16'h2C70 : rd_rsp_data <= 32'h00A8C754;
        16'h2C74 : rd_rsp_data <= 32'h0000C756;
        16'h2C80 : rd_rsp_data <= 32'h4C731AD5;
        16'h2C84 : rd_rsp_data <= 32'h3EE00000;
        16'h2C88 : rd_rsp_data <= 32'h005F7C00;
        16'h2C94 : rd_rsp_data <= 32'h00000050;
        16'h2C98 : rd_rsp_data <= 32'h08400000;
        16'h2CA8 : rd_rsp_data <= 32'h5E101006;
        16'h2CB0 : rd_rsp_data <= 32'h00004C64;
        16'h2CB4 : rd_rsp_data <= 32'h0000F7F3;
        16'h2CB8 : rd_rsp_data <= 32'h00002000;
        16'h2CC0 : rd_rsp_data <= 32'h000C0F0F;
        16'h2CC4 : rd_rsp_data <= 32'h301DB18F;
        16'h2CC8 : rd_rsp_data <= 32'h03CF0EB6;
        16'h2CCC : rd_rsp_data <= 32'h0056B814;
        16'h2CD0 : rd_rsp_data <= 32'h013C0980;
        16'h2CD4 : rd_rsp_data <= 32'hFBE7F77C;
        16'h2CD8 : rd_rsp_data <= 32'h2D495C3E;
        16'h2CDC : rd_rsp_data <= 32'h02A885DC;
        16'h2CE0 : rd_rsp_data <= 32'h028816A0;
        16'h2CE4 : rd_rsp_data <= 32'h02C2061D;
        16'h2CE8 : rd_rsp_data <= 32'h608060A6;
        16'h2CEC : rd_rsp_data <= 32'h007D7878;
        16'h2CF0 : rd_rsp_data <= 32'h31606060;
        16'h2CF4 : rd_rsp_data <= 32'h0062407F;
        16'h2CF8 : rd_rsp_data <= 32'h80313131;
        16'h2CFC : rd_rsp_data <= 32'h036060FF;
        16'h2D00 : rd_rsp_data <= 32'h00000001;
        16'h2D04 : rd_rsp_data <= 32'h000C3C3C;
        16'h2D0C : rd_rsp_data <= 32'h00000001;
        16'h2D10 : rd_rsp_data <= 32'h17171D1D;
        16'h2D1C : rd_rsp_data <= 32'h190F1622;
        16'h2D20 : rd_rsp_data <= 32'h052AAAD1;
        16'h2D80 : rd_rsp_data <= 32'h00000001;
        16'h2D84 : rd_rsp_data <= 32'h000C3C3C;
        16'h2D8C : rd_rsp_data <= 32'h00000001;
        16'h2D90 : rd_rsp_data <= 32'h17171D1D;
        16'h2D9C : rd_rsp_data <= 32'h190F1622;
        16'h2DA0 : rd_rsp_data <= 32'h052AAAD1;
        16'h2E00 : rd_rsp_data <= 32'h00000001;
        16'h2E04 : rd_rsp_data <= 32'h000C3C3C;
        16'h2E0C : rd_rsp_data <= 32'h00000001;
        16'h2E10 : rd_rsp_data <= 32'h17171D1D;
        16'h2E1C : rd_rsp_data <= 32'h190F1622;
        16'h2E20 : rd_rsp_data <= 32'h052AAAD1;
        16'h2E80 : rd_rsp_data <= 32'h00000001;
        16'h2E84 : rd_rsp_data <= 32'h000C3C3C;
        16'h2E8C : rd_rsp_data <= 32'h00000001;
        16'h2E90 : rd_rsp_data <= 32'h17171D1D;
        16'h2E9C : rd_rsp_data <= 32'h190F1622;
        16'h2EA0 : rd_rsp_data <= 32'h052AAAD1;
        16'h2F00 : rd_rsp_data <= 32'h00000001;
        16'h2F04 : rd_rsp_data <= 32'h000C3C3C;
        16'h2F0C : rd_rsp_data <= 32'h00000001;
        16'h2F10 : rd_rsp_data <= 32'h17171D1D;
        16'h2F1C : rd_rsp_data <= 32'h190F1622;
        16'h2F20 : rd_rsp_data <= 32'h052AAAD1;
        16'h2F80 : rd_rsp_data <= 32'h00000001;
        16'h2F84 : rd_rsp_data <= 32'h000C3C3C;
        16'h2F8C : rd_rsp_data <= 32'h00000001;
        16'h2F90 : rd_rsp_data <= 32'h17171D1D;
        16'h2F9C : rd_rsp_data <= 32'h190F1622;
        16'h2FA0 : rd_rsp_data <= 32'h052AAAD1;
        16'h3000 : rd_rsp_data <= 32'h00000001;
        16'h3004 : rd_rsp_data <= 32'h000C3C3C;
        16'h300C : rd_rsp_data <= 32'h00000001;
        16'h3010 : rd_rsp_data <= 32'h17171D1D;
        16'h301C : rd_rsp_data <= 32'h190F1622;
        16'h3020 : rd_rsp_data <= 32'h052AAAD1;
        16'h3080 : rd_rsp_data <= 32'h00000001;
        16'h3084 : rd_rsp_data <= 32'h000C3C3C;
        16'h308C : rd_rsp_data <= 32'h00000001;
        16'h3090 : rd_rsp_data <= 32'h17171D1D;
        16'h309C : rd_rsp_data <= 32'h190F1622;
        16'h30A0 : rd_rsp_data <= 32'h052AAAD1;
        16'h3100 : rd_rsp_data <= 32'h000C3C3C;
        16'h310C : rd_rsp_data <= 32'h00000001;
        16'h3110 : rd_rsp_data <= 32'h50000000;
        16'h3114 : rd_rsp_data <= 32'h60C02000;
        16'h3120 : rd_rsp_data <= 32'h08600080;
        16'h3124 : rd_rsp_data <= 32'h08600080;
        16'h3130 : rd_rsp_data <= 32'hE5B9FEF4;
        16'h3134 : rd_rsp_data <= 32'hF7B9FEF4;
        16'h3138 : rd_rsp_data <= 32'hE7FFC000;
        16'h313C : rd_rsp_data <= 32'h110F1622;
        16'h3140 : rd_rsp_data <= 32'h0B44A555;
        16'h3144 : rd_rsp_data <= 32'h007AC72B;
        16'h3148 : rd_rsp_data <= 32'h00000D3B;
        16'h3180 : rd_rsp_data <= 32'h000C3C3C;
        16'h318C : rd_rsp_data <= 32'h00000001;
        16'h3190 : rd_rsp_data <= 32'h50000000;
        16'h3194 : rd_rsp_data <= 32'h60C02000;
        16'h31A0 : rd_rsp_data <= 32'h08600080;
        16'h31A4 : rd_rsp_data <= 32'h08600080;
        16'h31B0 : rd_rsp_data <= 32'hDF77FCF4;
        16'h31B4 : rd_rsp_data <= 32'hE7FDDFE8;
        16'h31B8 : rd_rsp_data <= 32'hDFFDC000;
        16'h31BC : rd_rsp_data <= 32'h110F1622;
        16'h31C0 : rd_rsp_data <= 32'h0B44A555;
        16'h31C4 : rd_rsp_data <= 32'h007AC72B;
        16'h31C8 : rd_rsp_data <= 32'h00000D3B;
        16'h3200 : rd_rsp_data <= 32'h000C3C3C;
        16'h320C : rd_rsp_data <= 32'h00000001;
        16'h3210 : rd_rsp_data <= 32'h50000000;
        16'h3214 : rd_rsp_data <= 32'h60C02000;
        16'h3220 : rd_rsp_data <= 32'h08600080;
        16'h3224 : rd_rsp_data <= 32'h08600080;
        16'h3230 : rd_rsp_data <= 32'hE6B5FDE0;
        16'h3234 : rd_rsp_data <= 32'hFF3BBEFC;
        16'h3238 : rd_rsp_data <= 32'hFF7FE000;
        16'h323C : rd_rsp_data <= 32'h110F1622;
        16'h3240 : rd_rsp_data <= 32'h0B44A555;
        16'h3244 : rd_rsp_data <= 32'h007AC72B;
        16'h3248 : rd_rsp_data <= 32'h00000D3B;
        16'h3280 : rd_rsp_data <= 32'h000C3C3C;
        16'h328C : rd_rsp_data <= 32'h00000001;
        16'h3290 : rd_rsp_data <= 32'h50000000;
        16'h3294 : rd_rsp_data <= 32'h60C02000;
        16'h32A0 : rd_rsp_data <= 32'h08600080;
        16'h32A4 : rd_rsp_data <= 32'h08600080;
        16'h32B0 : rd_rsp_data <= 32'hFCF1DEF0;
        16'h32B4 : rd_rsp_data <= 32'hFF7DCE7C;
        16'h32B8 : rd_rsp_data <= 32'hE7F7B000;
        16'h32BC : rd_rsp_data <= 32'h110F1622;
        16'h32C0 : rd_rsp_data <= 32'h0B44A555;
        16'h32C4 : rd_rsp_data <= 32'h007AC72B;
        16'h32C8 : rd_rsp_data <= 32'h00000D3B;
        16'h3300 : rd_rsp_data <= 32'h28A00018;
        16'h3304 : rd_rsp_data <= 32'h70000221;
        16'h3308 : rd_rsp_data <= 32'h04003D2F;
        16'h3314 : rd_rsp_data <= 32'h18068682;
        16'h3318 : rd_rsp_data <= 32'h31E10013;
        16'h3320 : rd_rsp_data <= 32'h00000001;
        16'h3380 : rd_rsp_data <= 32'h00000001;
        16'h3384 : rd_rsp_data <= 32'h000C3C3C;
        16'h338C : rd_rsp_data <= 32'h00000001;
        16'h3390 : rd_rsp_data <= 32'h17171D1D;
        16'h339C : rd_rsp_data <= 32'h190F1622;
        16'h33A0 : rd_rsp_data <= 32'h052AAAD1;
        16'h3400 : rd_rsp_data <= 32'h00000001;
        16'h3404 : rd_rsp_data <= 32'h000C3C3C;
        16'h340C : rd_rsp_data <= 32'h00000001;
        16'h3410 : rd_rsp_data <= 32'h17171D1D;
        16'h341C : rd_rsp_data <= 32'h190F1622;
        16'h3420 : rd_rsp_data <= 32'h052AAAD1;
        16'h3480 : rd_rsp_data <= 32'h2001FC0B;
        16'h3484 : rd_rsp_data <= 32'h00000005;
        16'h3488 : rd_rsp_data <= 32'h009E0000;
        16'h348C : rd_rsp_data <= 32'h00800094;
        16'h3490 : rd_rsp_data <= 32'h00000100;
        16'h3494 : rd_rsp_data <= 32'h00000080;
        16'h3498 : rd_rsp_data <= 32'h057E4804;
        16'h349C : rd_rsp_data <= 32'h0000003B;
        16'h34A0 : rd_rsp_data <= 32'h8020E207;
        16'h34A4 : rd_rsp_data <= 32'h40155D63;
        16'h34A8 : rd_rsp_data <= 32'h00000075;
        16'h34AC : rd_rsp_data <= 32'h3FFE0000;
        16'h34B0 : rd_rsp_data <= 32'h0000020F;
        16'h34BC : rd_rsp_data <= 32'h60E7D545;
        16'h34C0 : rd_rsp_data <= 32'h0005C478;
        16'h34C8 : rd_rsp_data <= 32'h0E400010;
        16'h34D8 : rd_rsp_data <= 32'h0F000000;
        16'h34E0 : rd_rsp_data <= 32'h808D7887;
        16'h34E4 : rd_rsp_data <= 32'h7C89888C;
        16'h34E8 : rd_rsp_data <= 32'h78808D7C;
        16'h34EC : rd_rsp_data <= 32'hFF90857C;
        16'h34F0 : rd_rsp_data <= 32'h80808080;
        16'h34F4 : rd_rsp_data <= 32'h89852001;
        16'h3500 : rd_rsp_data <= 32'h00E20000;
        16'h3508 : rd_rsp_data <= 32'h00000006;
        16'h350C : rd_rsp_data <= 32'h0001CA00;
        16'h3510 : rd_rsp_data <= 32'h01660444;
        16'h3514 : rd_rsp_data <= 32'hE00DCE0C;
        16'h351C : rd_rsp_data <= 32'h08400000;
        16'h3534 : rd_rsp_data <= 32'h07500000;
        16'h3538 : rd_rsp_data <= 32'h82A885DC;
        16'h353C : rd_rsp_data <= 32'h028816A0;
        16'h3540 : rd_rsp_data <= 32'h02C2061D;
        16'h3544 : rd_rsp_data <= 32'h0154C222;
        16'h354C : rd_rsp_data <= 32'h01440000;
        16'h3550 : rd_rsp_data <= 32'hFFFF0000;
        16'h3554 : rd_rsp_data <= 32'h20000000;
        16'h3568 : rd_rsp_data <= 32'h000005EC;
        16'h357C : rd_rsp_data <= 32'h00062000;
        16'h3580 : rd_rsp_data <= 32'h2001FC0B;
        16'h3584 : rd_rsp_data <= 32'h00000005;
        16'h3588 : rd_rsp_data <= 32'h009C0000;
        16'h358C : rd_rsp_data <= 32'h00800092;
        16'h3590 : rd_rsp_data <= 32'h00000100;
        16'h3594 : rd_rsp_data <= 32'h00000080;
        16'h3598 : rd_rsp_data <= 32'h057E4804;
        16'h359C : rd_rsp_data <= 32'h0000003B;
        16'h35A0 : rd_rsp_data <= 32'h8020F207;
        16'h35A4 : rd_rsp_data <= 32'h40155D63;
        16'h35A8 : rd_rsp_data <= 32'h00000075;
        16'h35AC : rd_rsp_data <= 32'h3FFE0000;
        16'h35B0 : rd_rsp_data <= 32'h0000020F;
        16'h35BC : rd_rsp_data <= 32'h60E7D545;
        16'h35C0 : rd_rsp_data <= 32'h0005C478;
        16'h35C8 : rd_rsp_data <= 32'h0E400010;
        16'h35D8 : rd_rsp_data <= 32'h0F000000;
        16'h35E0 : rd_rsp_data <= 32'h808F8887;
        16'h35E4 : rd_rsp_data <= 32'h9B918F7C;
        16'h35E8 : rd_rsp_data <= 32'h8B89918B;
        16'h35EC : rd_rsp_data <= 32'hFF94899C;
        16'h35F0 : rd_rsp_data <= 32'h80808080;
        16'h35F4 : rd_rsp_data <= 32'h98902001;
        16'h3600 : rd_rsp_data <= 32'h00E20000;
        16'h3608 : rd_rsp_data <= 32'h00000006;
        16'h360C : rd_rsp_data <= 32'h0001CA00;
        16'h3610 : rd_rsp_data <= 32'h01660444;
        16'h3614 : rd_rsp_data <= 32'hE00DCE0C;
        16'h361C : rd_rsp_data <= 32'h08400000;
        16'h3634 : rd_rsp_data <= 32'h07500000;
        16'h3638 : rd_rsp_data <= 32'h82A885DC;
        16'h363C : rd_rsp_data <= 32'h028816A0;
        16'h3640 : rd_rsp_data <= 32'h02C2061D;
        16'h3644 : rd_rsp_data <= 32'h0154C222;
        16'h364C : rd_rsp_data <= 32'h01440000;
        16'h3650 : rd_rsp_data <= 32'hFFFF0000;
        16'h3654 : rd_rsp_data <= 32'h20000000;
        16'h367C : rd_rsp_data <= 32'h00062000;
        16'h3680 : rd_rsp_data <= 32'h2001A07F;
        16'h3684 : rd_rsp_data <= 32'h00000005;
        16'h3688 : rd_rsp_data <= 32'h00900000;
        16'h368C : rd_rsp_data <= 32'h00000080;
        16'h3690 : rd_rsp_data <= 32'h00000100;
        16'h3698 : rd_rsp_data <= 32'h057E4804;
        16'h369C : rd_rsp_data <= 32'h0000003B;
        16'h36A0 : rd_rsp_data <= 32'h8020F207;
        16'h36A4 : rd_rsp_data <= 32'h40155D63;
        16'h36A8 : rd_rsp_data <= 32'h00000075;
        16'h36AC : rd_rsp_data <= 32'h3FFE0000;
        16'h36B0 : rd_rsp_data <= 32'h0000020F;
        16'h36BC : rd_rsp_data <= 32'h60E7D545;
        16'h36C0 : rd_rsp_data <= 32'h0005C478;
        16'h36C8 : rd_rsp_data <= 32'h0E400010;
        16'h36D8 : rd_rsp_data <= 32'h0F000000;
        16'h36E0 : rd_rsp_data <= 32'h80949878;
        16'h36E4 : rd_rsp_data <= 32'h85889C93;
        16'h36E8 : rd_rsp_data <= 32'h8E8D917C;
        16'h36EC : rd_rsp_data <= 32'hFF97889F;
        16'h36F0 : rd_rsp_data <= 32'h80808080;
        16'h36F4 : rd_rsp_data <= 32'h8D8C2001;
        16'h3700 : rd_rsp_data <= 32'h00E20000;
        16'h3708 : rd_rsp_data <= 32'h00000006;
        16'h370C : rd_rsp_data <= 32'h0001CA00;
        16'h3710 : rd_rsp_data <= 32'h01660444;
        16'h3714 : rd_rsp_data <= 32'hE00DCE0C;
        16'h371C : rd_rsp_data <= 32'h08400000;
        16'h3734 : rd_rsp_data <= 32'h07500000;
        16'h3738 : rd_rsp_data <= 32'h82A885DC;
        16'h373C : rd_rsp_data <= 32'h028816A0;
        16'h3740 : rd_rsp_data <= 32'h02C2061D;
        16'h3744 : rd_rsp_data <= 32'h0154C222;
        16'h374C : rd_rsp_data <= 32'h01440000;
        16'h3750 : rd_rsp_data <= 32'hFFFF0000;
        16'h3754 : rd_rsp_data <= 32'h20000000;
        16'h3768 : rd_rsp_data <= 32'h00000526;
        16'h377C : rd_rsp_data <= 32'h00062000;
        16'h3780 : rd_rsp_data <= 32'h2001A07F;
        16'h3784 : rd_rsp_data <= 32'h00000005;
        16'h3788 : rd_rsp_data <= 32'h00880000;
        16'h378C : rd_rsp_data <= 32'h00000080;
        16'h3790 : rd_rsp_data <= 32'h00000100;
        16'h3798 : rd_rsp_data <= 32'h057E4804;
        16'h379C : rd_rsp_data <= 32'h0000003B;
        16'h37A0 : rd_rsp_data <= 32'h8020E207;
        16'h37A4 : rd_rsp_data <= 32'h40155D63;
        16'h37A8 : rd_rsp_data <= 32'h00000075;
        16'h37AC : rd_rsp_data <= 32'h3FFE0000;
        16'h37B0 : rd_rsp_data <= 32'h0000020F;
        16'h37BC : rd_rsp_data <= 32'h60E7D545;
        16'h37C0 : rd_rsp_data <= 32'h0005C478;
        16'h37C8 : rd_rsp_data <= 32'h0E400010;
        16'h37D8 : rd_rsp_data <= 32'h0F000000;
        16'h37E0 : rd_rsp_data <= 32'h808D877C;
        16'h37E4 : rd_rsp_data <= 32'h898C9489;
        16'h37E8 : rd_rsp_data <= 32'h907E7C78;
        16'h37EC : rd_rsp_data <= 32'hFF98808D;
        16'h37F0 : rd_rsp_data <= 32'h80808080;
        16'h37F4 : rd_rsp_data <= 32'h8F942001;
        16'h3800 : rd_rsp_data <= 32'h00E20000;
        16'h380C : rd_rsp_data <= 32'h0001CA00;
        16'h3810 : rd_rsp_data <= 32'h01660444;
        16'h3814 : rd_rsp_data <= 32'hE00DCE0C;
        16'h381C : rd_rsp_data <= 32'h08400000;
        16'h3834 : rd_rsp_data <= 32'h07500000;
        16'h3838 : rd_rsp_data <= 32'h82A885DC;
        16'h383C : rd_rsp_data <= 32'h028816A0;
        16'h3840 : rd_rsp_data <= 32'h02C2061D;
        16'h3844 : rd_rsp_data <= 32'h0154C222;
        16'h384C : rd_rsp_data <= 32'h01440000;
        16'h3850 : rd_rsp_data <= 32'hFFFF0000;
        16'h3854 : rd_rsp_data <= 32'h20000000;
        16'h3868 : rd_rsp_data <= 32'h0000069E;
        16'h387C : rd_rsp_data <= 32'h00002000;
        16'h3880 : rd_rsp_data <= 32'h2001F590;
        16'h3884 : rd_rsp_data <= 32'h00000005;
        16'h3888 : rd_rsp_data <= 32'h007E0000;
        16'h388C : rd_rsp_data <= 32'h00800080;
        16'h3890 : rd_rsp_data <= 32'h00000100;
        16'h3898 : rd_rsp_data <= 32'h057E4804;
        16'h389C : rd_rsp_data <= 32'h0000003B;
        16'h38A0 : rd_rsp_data <= 32'h8020E607;
        16'h38A4 : rd_rsp_data <= 32'h40155D63;
        16'h38A8 : rd_rsp_data <= 32'h00000075;
        16'h38AC : rd_rsp_data <= 32'h3FFE0000;
        16'h38B0 : rd_rsp_data <= 32'h0000020F;
        16'h38BC : rd_rsp_data <= 32'h60E7D545;
        16'h38C0 : rd_rsp_data <= 32'h0005C478;
        16'h38C8 : rd_rsp_data <= 32'h0E400010;
        16'h38D8 : rd_rsp_data <= 32'h0F000000;
        16'h38E0 : rd_rsp_data <= 32'h80928F68;
        16'h38E4 : rd_rsp_data <= 32'h87909094;
        16'h38E8 : rd_rsp_data <= 32'h89878185;
        16'h38EC : rd_rsp_data <= 32'hFF909089;
        16'h38F0 : rd_rsp_data <= 32'h80808080;
        16'h38F4 : rd_rsp_data <= 32'h7C802001;
        16'h3900 : rd_rsp_data <= 32'h00E20000;
        16'h3908 : rd_rsp_data <= 32'h00000006;
        16'h390C : rd_rsp_data <= 32'h0001CA00;
        16'h3910 : rd_rsp_data <= 32'h01660444;
        16'h3914 : rd_rsp_data <= 32'hE00DCE0C;
        16'h391C : rd_rsp_data <= 32'h08400000;
        16'h3934 : rd_rsp_data <= 32'h07500000;
        16'h3938 : rd_rsp_data <= 32'h82A885DC;
        16'h393C : rd_rsp_data <= 32'h028816A0;
        16'h3940 : rd_rsp_data <= 32'h02C2061D;
        16'h3944 : rd_rsp_data <= 32'h0154C222;
        16'h394C : rd_rsp_data <= 32'h01440000;
        16'h3950 : rd_rsp_data <= 32'hFFFF0000;
        16'h3954 : rd_rsp_data <= 32'h20000000;
        16'h3968 : rd_rsp_data <= 32'h0000037C;
        16'h397C : rd_rsp_data <= 32'h00062000;
        16'h3980 : rd_rsp_data <= 32'h2001F470;
        16'h3984 : rd_rsp_data <= 32'h00000005;
        16'h3988 : rd_rsp_data <= 32'h00820000;
        16'h398C : rd_rsp_data <= 32'h00800080;
        16'h3990 : rd_rsp_data <= 32'h00000100;
        16'h3998 : rd_rsp_data <= 32'h057E4804;
        16'h399C : rd_rsp_data <= 32'h0000003B;
        16'h39A0 : rd_rsp_data <= 32'h8020F207;
        16'h39A4 : rd_rsp_data <= 32'h40155D63;
        16'h39A8 : rd_rsp_data <= 32'h00000075;
        16'h39AC : rd_rsp_data <= 32'h3FFE0000;
        16'h39B0 : rd_rsp_data <= 32'h0000020F;
        16'h39BC : rd_rsp_data <= 32'h60E7D545;
        16'h39C0 : rd_rsp_data <= 32'h0005C478;
        16'h39C8 : rd_rsp_data <= 32'h0E400010;
        16'h39D8 : rd_rsp_data <= 32'h0F000000;
        16'h39E0 : rd_rsp_data <= 32'h80939478;
        16'h39E4 : rd_rsp_data <= 32'h7C9C918F;
        16'h39E8 : rd_rsp_data <= 32'h9885857E;
        16'h39EC : rd_rsp_data <= 32'hFF94919F;
        16'h39F0 : rd_rsp_data <= 32'h80808080;
        16'h39F4 : rd_rsp_data <= 32'h93982001;
        16'h3A00 : rd_rsp_data <= 32'h00E20000;
        16'h3A0C : rd_rsp_data <= 32'h0001CA00;
        16'h3A10 : rd_rsp_data <= 32'h01660444;
        16'h3A14 : rd_rsp_data <= 32'hE00DCE0C;
        16'h3A1C : rd_rsp_data <= 32'h08400000;
        16'h3A34 : rd_rsp_data <= 32'h07500000;
        16'h3A38 : rd_rsp_data <= 32'h82A885DC;
        16'h3A3C : rd_rsp_data <= 32'h028816A0;
        16'h3A40 : rd_rsp_data <= 32'h02C2061D;
        16'h3A44 : rd_rsp_data <= 32'h0154C222;
        16'h3A4C : rd_rsp_data <= 32'h01440000;
        16'h3A50 : rd_rsp_data <= 32'hFFFF0000;
        16'h3A54 : rd_rsp_data <= 32'h20000000;
        16'h3A7C : rd_rsp_data <= 32'h00002000;
        16'h3A80 : rd_rsp_data <= 32'h2001D61F;
        16'h3A84 : rd_rsp_data <= 32'h00000005;
        16'h3A88 : rd_rsp_data <= 32'h00920000;
        16'h3A8C : rd_rsp_data <= 32'h00880080;
        16'h3A90 : rd_rsp_data <= 32'h00000100;
        16'h3A98 : rd_rsp_data <= 32'h057E4804;
        16'h3A9C : rd_rsp_data <= 32'h0000003B;
        16'h3AA0 : rd_rsp_data <= 32'h8020E607;
        16'h3AA4 : rd_rsp_data <= 32'h40155D63;
        16'h3AA8 : rd_rsp_data <= 32'h00000075;
        16'h3AAC : rd_rsp_data <= 32'h3FFE0000;
        16'h3AB0 : rd_rsp_data <= 32'h0000020F;
        16'h3ABC : rd_rsp_data <= 32'h60E7D545;
        16'h3AC0 : rd_rsp_data <= 32'h0005C478;
        16'h3AC8 : rd_rsp_data <= 32'h0E400010;
        16'h3AD8 : rd_rsp_data <= 32'h0F000000;
        16'h3AE0 : rd_rsp_data <= 32'h80939079;
        16'h3AE4 : rd_rsp_data <= 32'h7C939889;
        16'h3AE8 : rd_rsp_data <= 32'hA0787E8F;
        16'h3AEC : rd_rsp_data <= 32'hFFA07888;
        16'h3AF0 : rd_rsp_data <= 32'h80808080;
        16'h3AF4 : rd_rsp_data <= 32'h8B7C2001;
        16'h3B00 : rd_rsp_data <= 32'h00E20000;
        16'h3B08 : rd_rsp_data <= 32'h00000002;
        16'h3B0C : rd_rsp_data <= 32'h0001CA00;
        16'h3B10 : rd_rsp_data <= 32'h01660444;
        16'h3B14 : rd_rsp_data <= 32'hE00DCE0C;
        16'h3B1C : rd_rsp_data <= 32'h08400000;
        16'h3B34 : rd_rsp_data <= 32'h07500000;
        16'h3B38 : rd_rsp_data <= 32'h82A885DC;
        16'h3B3C : rd_rsp_data <= 32'h028816A0;
        16'h3B40 : rd_rsp_data <= 32'h02C2061D;
        16'h3B44 : rd_rsp_data <= 32'h0154C222;
        16'h3B4C : rd_rsp_data <= 32'h01440000;
        16'h3B50 : rd_rsp_data <= 32'hFFFF0000;
        16'h3B54 : rd_rsp_data <= 32'h20000000;
        16'h3B68 : rd_rsp_data <= 32'h00000554;
        16'h3B7C : rd_rsp_data <= 32'h00022000;
        16'h3B80 : rd_rsp_data <= 32'h2001D61F;
        16'h3B84 : rd_rsp_data <= 32'h00000005;
        16'h3B88 : rd_rsp_data <= 32'h00860000;
        16'h3B8C : rd_rsp_data <= 32'h00940080;
        16'h3B90 : rd_rsp_data <= 32'h00000100;
        16'h3B98 : rd_rsp_data <= 32'h057E4804;
        16'h3B9C : rd_rsp_data <= 32'h0000003B;
        16'h3BA0 : rd_rsp_data <= 32'h8020E607;
        16'h3BA4 : rd_rsp_data <= 32'h40155D63;
        16'h3BA8 : rd_rsp_data <= 32'h00000075;
        16'h3BAC : rd_rsp_data <= 32'h3FFE0000;
        16'h3BB0 : rd_rsp_data <= 32'h0000020F;
        16'h3BBC : rd_rsp_data <= 32'h60E7D545;
        16'h3BC0 : rd_rsp_data <= 32'h0005C478;
        16'h3BC8 : rd_rsp_data <= 32'h0E400010;
        16'h3BD8 : rd_rsp_data <= 32'h0F000000;
        16'h3BE0 : rd_rsp_data <= 32'h80937C89;
        16'h3BE4 : rd_rsp_data <= 32'h95989894;
        16'h3BE8 : rd_rsp_data <= 32'h87898593;
        16'h3BEC : rd_rsp_data <= 32'hFF8C9090;
        16'h3BF0 : rd_rsp_data <= 32'h80808080;
        16'h3BF4 : rd_rsp_data <= 32'h888D2001;
        16'h3C00 : rd_rsp_data <= 32'h00E20000;
        16'h3C08 : rd_rsp_data <= 32'h00000004;
        16'h3C0C : rd_rsp_data <= 32'h0001CA00;
        16'h3C10 : rd_rsp_data <= 32'h01660444;
        16'h3C14 : rd_rsp_data <= 32'hE00DCE0C;
        16'h3C1C : rd_rsp_data <= 32'h08400000;
        16'h3C34 : rd_rsp_data <= 32'h07500000;
        16'h3C38 : rd_rsp_data <= 32'h82A885DC;
        16'h3C3C : rd_rsp_data <= 32'h028816A0;
        16'h3C40 : rd_rsp_data <= 32'h02C2061D;
        16'h3C44 : rd_rsp_data <= 32'h0154C222;
        16'h3C4C : rd_rsp_data <= 32'h01440000;
        16'h3C50 : rd_rsp_data <= 32'hFFFF0000;
        16'h3C54 : rd_rsp_data <= 32'h20000000;
        16'h3C68 : rd_rsp_data <= 32'h00000662;
        16'h3C7C : rd_rsp_data <= 32'h00042000;
        16'h3C80 : rd_rsp_data <= 32'h78444842;
        16'h3C84 : rd_rsp_data <= 32'h05800035;
        16'h3C88 : rd_rsp_data <= 32'h17171D1D;
        16'h3C8C : rd_rsp_data <= 32'h0154C222;
        16'h3C90 : rd_rsp_data <= 32'h00004229;
        16'h3C94 : rd_rsp_data <= 32'h20480000;
        16'h3C9C : rd_rsp_data <= 32'h007C201E;
        16'h3CA0 : rd_rsp_data <= 32'h2C2C2C2C;
        16'h3CA4 : rd_rsp_data <= 32'h00042C2C;
        16'h3CBC : rd_rsp_data <= 32'h00000001;
        16'h3CD4 : rd_rsp_data <= 32'h00008080;
        16'h3CE8 : rd_rsp_data <= 32'h00000103;
        16'h3CF0 : rd_rsp_data <= 32'h03DF7B01;
        16'h3D00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3D9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3DFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h3E00 : rd_rsp_data <= 32'h003E0F1D;
        16'h3E04 : rd_rsp_data <= 32'h003E0F1D;
        16'h3E08 : rd_rsp_data <= 32'h003E0F1D;
        16'h3E0C : rd_rsp_data <= 32'h003E0F1D;
        16'h3E10 : rd_rsp_data <= 32'h003E0F1D;
        16'h3E14 : rd_rsp_data <= 32'h003E0F1D;
        16'h3E18 : rd_rsp_data <= 32'h003E0F1D;
        16'h3E1C : rd_rsp_data <= 32'h003E0F1D;
        16'h3E20 : rd_rsp_data <= 32'h00000200;
        16'h3E24 : rd_rsp_data <= 32'h7C64217A;
        16'h3E28 : rd_rsp_data <= 32'hE1642130;
        16'h3E2C : rd_rsp_data <= 32'h7FE00D9F;
        16'h3E30 : rd_rsp_data <= 32'h7FE00D9F;
        16'h3E34 : rd_rsp_data <= 32'h7FE00C9D;
        16'h3E38 : rd_rsp_data <= 32'h7FE00C9D;
        16'h3E3C : rd_rsp_data <= 32'h7FE00D9F;
        16'h3E40 : rd_rsp_data <= 32'h7FE00D9F;
        16'h3E44 : rd_rsp_data <= 32'h7FE00C9D;
        16'h3E48 : rd_rsp_data <= 32'h7FE00C9D;
        16'h3E4C : rd_rsp_data <= 32'h4561E000;
        16'h3E50 : rd_rsp_data <= 32'h4561E000;
        16'h3E54 : rd_rsp_data <= 32'h4539C000;
        16'h3E58 : rd_rsp_data <= 32'h4539C000;
        16'h3E5C : rd_rsp_data <= 32'h4561F000;
        16'h3E60 : rd_rsp_data <= 32'h4561F000;
        16'h3E64 : rd_rsp_data <= 32'h4539D000;
        16'h3E68 : rd_rsp_data <= 32'h4539D000;
        16'h3EA0 : rd_rsp_data <= 32'h00000908;
        16'h3EC4 : rd_rsp_data <= 32'h00000400;
        16'h3EC8 : rd_rsp_data <= 32'h00000001;
        16'h3ECC : rd_rsp_data <= 32'h000004E4;
        16'h3ED4 : rd_rsp_data <= 32'h00000001;
        16'h3ED8 : rd_rsp_data <= 32'h47200000;
        16'h3F80 : rd_rsp_data <= 32'h01000208;
        16'h3F84 : rd_rsp_data <= 32'h00000400;
        16'h3F88 : rd_rsp_data <= 32'h0100060A;
        16'h3F8C : rd_rsp_data <= 32'h00000400;
        16'h4000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h400C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h401C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h402C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h403C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h404C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h405C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h406C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h407C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h408C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h409C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h40FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h410C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h411C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h412C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h413C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h414C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h415C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h416C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h417C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h418C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h419C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h41FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h420C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h421C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h422C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h423C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h424C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h425C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h426C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h427C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h428C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h429C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h42FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h430C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h431C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h432C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h433C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h434C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h435C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h436C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h437C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h438C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h439C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h43FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h440C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h441C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h442C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h443C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h444C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h445C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h446C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h447C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h448C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h449C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h44FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h450C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h451C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h452C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h453C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h454C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h455C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h456C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h457C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h458C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h459C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h45FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h460C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h461C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h462C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h463C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h464C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h465C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h466C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h467C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h468C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h469C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h46FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h470C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h471C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h472C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h473C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h474C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h475C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h476C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h477C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h478C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h479C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h47FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h480C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h481C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h482C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h483C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h484C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h485C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h486C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h487C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h488C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h489C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h48FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h490C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h491C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h492C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h493C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h494C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h495C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h496C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h497C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h498C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h499C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h49FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4A9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4ABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4ACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4ADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4AFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4B9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4BFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4C9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4CFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4D9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4DFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4E9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4ECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4ED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4ED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4ED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4EFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4F9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h4FFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h500C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h501C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h502C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h503C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h504C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h505C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h506C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h507C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h508C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h509C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h50FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h510C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h511C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h512C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h513C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h514C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h515C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h516C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h517C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h518C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h519C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h51FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h520C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h521C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h522C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h523C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h524C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h525C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h526C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h527C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h528C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h529C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h52FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h530C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h531C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h532C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h533C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h534C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h535C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h536C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h537C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h538C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h539C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h53FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5400 : rd_rsp_data <= 32'hFED90001;
        16'h5410 : rd_rsp_data <= 32'hFED91001;
        16'h5418 : rd_rsp_data <= 32'h00000010;
        16'h541C : rd_rsp_data <= 32'h30000000;
        16'h5428 : rd_rsp_data <= 32'h00000004;
        16'h54A0 : rd_rsp_data <= 32'h03102001;
        16'h5520 : rd_rsp_data <= 32'h01000208;
        16'h5524 : rd_rsp_data <= 32'h00000400;
        16'h5528 : rd_rsp_data <= 32'h0100820A;
        16'h552C : rd_rsp_data <= 32'h00000408;
        16'h5530 : rd_rsp_data <= 32'h0100820A;
        16'h5534 : rd_rsp_data <= 32'h00000408;
        16'h5538 : rd_rsp_data <= 32'h01000200;
        16'h553C : rd_rsp_data <= 32'h00000400;
        16'h5548 : rd_rsp_data <= 32'h01000200;
        16'h554C : rd_rsp_data <= 32'h00000400;
        16'h5550 : rd_rsp_data <= 32'h01010208;
        16'h5554 : rd_rsp_data <= 32'h00000400;
        16'h5560 : rd_rsp_data <= 32'h0101821F;
        16'h5564 : rd_rsp_data <= 32'h00001C08;
        16'h5568 : rd_rsp_data <= 32'h01000208;
        16'h556C : rd_rsp_data <= 32'h00000400;
        16'h5570 : rd_rsp_data <= 32'h00000400;
        16'h5578 : rd_rsp_data <= 32'h01000208;
        16'h557C : rd_rsp_data <= 32'h00000400;
        16'h5580 : rd_rsp_data <= 32'h01008208;
        16'h5584 : rd_rsp_data <= 32'h00000408;
        16'h5588 : rd_rsp_data <= 32'h01008208;
        16'h558C : rd_rsp_data <= 32'h00000408;
        16'h5590 : rd_rsp_data <= 32'h01000208;
        16'h5594 : rd_rsp_data <= 32'h00000400;
        16'h5598 : rd_rsp_data <= 32'h0100021A;
        16'h559C : rd_rsp_data <= 32'h00000400;
        16'h5824 : rd_rsp_data <= 32'h00000055;
        16'h5828 : rd_rsp_data <= 32'h47CE7C61;
        16'h582C : rd_rsp_data <= 32'h0000007C;
        16'h5830 : rd_rsp_data <= 32'h36CD9CF3;
        16'h5834 : rd_rsp_data <= 32'h00000032;
        16'h5838 : rd_rsp_data <= 32'h0000EA18;
        16'h5840 : rd_rsp_data <= 32'h0000EA18;
        16'h5848 : rd_rsp_data <= 32'h00009E66;
        16'h5850 : rd_rsp_data <= 32'h00009E66;
        16'h5858 : rd_rsp_data <= 32'h00005561;
        16'h5860 : rd_rsp_data <= 32'h39963250;
        16'h5864 : rd_rsp_data <= 32'h0000070B;
        16'h5868 : rd_rsp_data <= 32'h0009B274;
        16'h5870 : rd_rsp_data <= 32'h00066D6E;
        16'h5880 : rd_rsp_data <= 32'h00000040;
        16'h588C : rd_rsp_data <= 32'h00000001;
        16'h58A4 : rd_rsp_data <= 32'h00000002;
        16'h58A8 : rd_rsp_data <= 32'h00001327;
        16'h58FC : rd_rsp_data <= 32'h18021000;
        16'h5904 : rd_rsp_data <= 32'h01020000;
        16'h5918 : rd_rsp_data <= 32'h27000463;
        16'h591C : rd_rsp_data <= 32'h001A1B20;
        16'h5920 : rd_rsp_data <= 32'h00000010;
        16'h5924 : rd_rsp_data <= 32'h00000010;
        16'h5928 : rd_rsp_data <= 32'h204F1068;
        16'h592C : rd_rsp_data <= 32'h00000011;
        16'h5930 : rd_rsp_data <= 32'h000001B8;
        16'h5938 : rd_rsp_data <= 32'h000A0E03;
        16'h593C : rd_rsp_data <= 32'h54B10200;
        16'h5954 : rd_rsp_data <= 32'h00040000;
        16'h5958 : rd_rsp_data <= 32'hF1811C00;
        16'h595C : rd_rsp_data <= 32'h0004083D;
        16'h5968 : rd_rsp_data <= 32'h93501839;
        16'h596C : rd_rsp_data <= 32'h0FC04D29;
        16'h5974 : rd_rsp_data <= 32'h0000EA18;
        16'h5984 : rd_rsp_data <= 32'hE2ACD64B;
        16'h5994 : rd_rsp_data <= 32'h000000FF;
        16'h5998 : rd_rsp_data <= 32'h0006061F;
        16'h59A0 : rd_rsp_data <= 32'h00DF8370;
        16'h59A4 : rd_rsp_data <= 32'h004283C0;
        16'h59C0 : rd_rsp_data <= 32'h881E0000;
        16'h59D0 : rd_rsp_data <= 32'h1737691E;
        16'h59D4 : rd_rsp_data <= 32'h000009EF;
        16'h59D8 : rd_rsp_data <= 32'h529757F9;
        16'h59DC : rd_rsp_data <= 32'h00000059;
        16'h59E0 : rd_rsp_data <= 32'h59EF028E;
        16'h59E4 : rd_rsp_data <= 32'h00000059;
        16'h59E8 : rd_rsp_data <= 32'h7F56A1F0;
        16'h59EC : rd_rsp_data <= 32'h000006F7;
        16'h59F0 : rd_rsp_data <= 32'h0009E660;
        16'h59F8 : rd_rsp_data <= 32'h00005561;
        16'h5A08 : rd_rsp_data <= 32'h00000108;
        16'h5A0C : rd_rsp_data <= 32'h00333312;
        16'h5A10 : rd_rsp_data <= 32'h000001D3;
        16'h5A14 : rd_rsp_data <= 32'h00113004;
        16'h5A18 : rd_rsp_data <= 32'h003A0A33;
        16'h5A28 : rd_rsp_data <= 32'h6D92434B;
        16'h5A2C : rd_rsp_data <= 32'h00000059;
        16'h5A30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5A34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5A38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5B04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h5B10 : rd_rsp_data <= 32'h800000FF;
        16'h5C14 : rd_rsp_data <= 32'h00003008;
        16'h5C18 : rd_rsp_data <= 32'h00000610;
        16'h5C30 : rd_rsp_data <= 32'h27000463;
        16'h5C34 : rd_rsp_data <= 32'h001A1B20;
        16'h5D10 : rd_rsp_data <= 32'h00000002;
        16'h5D20 : rd_rsp_data <= 32'h00000005;
        16'h5D24 : rd_rsp_data <= 32'h000001F4;
        16'h5D34 : rd_rsp_data <= 32'h881E881E;
        16'h5D38 : rd_rsp_data <= 32'h881E881E;
        16'h5D48 : rd_rsp_data <= 32'h00011000;
        16'h5D54 : rd_rsp_data <= 32'h00000011;
        16'h5D60 : rd_rsp_data <= 32'h00000100;
        16'h5D70 : rd_rsp_data <= 32'h49400000;
        16'h5D78 : rd_rsp_data <= 32'h00000001;
        16'h5D7C : rd_rsp_data <= 32'h00004000;
        16'h5DA0 : rd_rsp_data <= 32'h0000006C;
        16'h5DA8 : rd_rsp_data <= 32'h00000003;
        16'h5DB0 : rd_rsp_data <= 32'h49400000;
        16'h5DB8 : rd_rsp_data <= 32'h00000001;
        16'h5DBC : rd_rsp_data <= 32'h00008000;
        16'h5DD0 : rd_rsp_data <= 32'h49407000;
        16'h5DD8 : rd_rsp_data <= 32'h00000006;
        16'h5DDC : rd_rsp_data <= 32'h00000034;
        16'h5E00 : rd_rsp_data <= 32'h39B81118;
        16'h5E04 : rd_rsp_data <= 32'h39B81118;
        16'h5EF0 : rd_rsp_data <= 32'h1F000600;
        16'h5F00 : rd_rsp_data <= 32'h00002106;
        16'h5F04 : rd_rsp_data <= 32'h00000011;
        16'h5F08 : rd_rsp_data <= 32'h00000014;
        16'h5F18 : rd_rsp_data <= 32'h00000001;
        16'h5F3C : rd_rsp_data <= 32'h0000001A;
        16'h5F40 : rd_rsp_data <= 32'h00160168;
        16'h5F48 : rd_rsp_data <= 32'h001C0208;
        16'h5F54 : rd_rsp_data <= 32'h00000019;
        16'h5F60 : rd_rsp_data <= 32'h000185AC;
        16'h5F70 : rd_rsp_data <= 32'h00000001;
        16'h5F74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6000 : rd_rsp_data <= 32'h00000044;
        16'h6004 : rd_rsp_data <= 32'h8000007F;
        16'h6008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6040 : rd_rsp_data <= 32'h130C3200;
        16'h6048 : rd_rsp_data <= 32'h00008001;
        16'h604C : rd_rsp_data <= 32'h00000100;
        16'h6050 : rd_rsp_data <= 32'h00000100;
        16'h6054 : rd_rsp_data <= 32'h10000800;
        16'h6058 : rd_rsp_data <= 32'h10000800;
        16'h605C : rd_rsp_data <= 32'h00000001;
        16'h61B0 : rd_rsp_data <= 32'h130C3200;
        16'h61B8 : rd_rsp_data <= 32'h00008001;
        16'h61BC : rd_rsp_data <= 32'h00000100;
        16'h61C0 : rd_rsp_data <= 32'h00000100;
        16'h61C4 : rd_rsp_data <= 32'h10000800;
        16'h61C8 : rd_rsp_data <= 32'h10000800;
        16'h61CC : rd_rsp_data <= 32'h13082400;
        16'h61D0 : rd_rsp_data <= 32'h00010000;
        16'h6200 : rd_rsp_data <= 32'h00000044;
        16'h6204 : rd_rsp_data <= 32'h8000007F;
        16'h6208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6240 : rd_rsp_data <= 32'h130C3200;
        16'h6248 : rd_rsp_data <= 32'h00008001;
        16'h624C : rd_rsp_data <= 32'h00000100;
        16'h6250 : rd_rsp_data <= 32'h00000100;
        16'h6254 : rd_rsp_data <= 32'h10000800;
        16'h6258 : rd_rsp_data <= 32'h10000800;
        16'h625C : rd_rsp_data <= 32'h00000001;
        16'h63B0 : rd_rsp_data <= 32'h130C3200;
        16'h63B8 : rd_rsp_data <= 32'h00008001;
        16'h63BC : rd_rsp_data <= 32'h00000100;
        16'h63C0 : rd_rsp_data <= 32'h00000100;
        16'h63C4 : rd_rsp_data <= 32'h10000800;
        16'h63C8 : rd_rsp_data <= 32'h10000800;
        16'h63CC : rd_rsp_data <= 32'h13082400;
        16'h63D0 : rd_rsp_data <= 32'h00010000;
        16'h6800 : rd_rsp_data <= 32'h01000208;
        16'h6804 : rd_rsp_data <= 32'h00000400;
        16'h6808 : rd_rsp_data <= 32'h0100020A;
        16'h680C : rd_rsp_data <= 32'h00000400;
        16'h6810 : rd_rsp_data <= 32'h0100020A;
        16'h6814 : rd_rsp_data <= 32'h00000400;
        16'h6818 : rd_rsp_data <= 32'h01000208;
        16'h681C : rd_rsp_data <= 32'h00000400;
        16'h6820 : rd_rsp_data <= 32'h00000400;
        16'h6828 : rd_rsp_data <= 32'h01000208;
        16'h682C : rd_rsp_data <= 32'h00000400;
        16'h6830 : rd_rsp_data <= 32'h0100021A;
        16'h6834 : rd_rsp_data <= 32'h00000400;
        16'h6850 : rd_rsp_data <= 32'h0100020A;
        16'h6854 : rd_rsp_data <= 32'h00000400;
        16'h6858 : rd_rsp_data <= 32'h0100020A;
        16'h685C : rd_rsp_data <= 32'h00000400;
        16'h6860 : rd_rsp_data <= 32'h0100020A;
        16'h6864 : rd_rsp_data <= 32'h00000400;
        16'h6878 : rd_rsp_data <= 32'h0100020A;
        16'h687C : rd_rsp_data <= 32'h00000400;
        16'h6880 : rd_rsp_data <= 32'h0100020A;
        16'h6884 : rd_rsp_data <= 32'h00000400;
        16'h6888 : rd_rsp_data <= 32'h0100020A;
        16'h688C : rd_rsp_data <= 32'h00000400;
        16'h6890 : rd_rsp_data <= 32'h01000208;
        16'h6894 : rd_rsp_data <= 32'h00000400;
        16'h6898 : rd_rsp_data <= 32'h0100020A;
        16'h689C : rd_rsp_data <= 32'h00000400;
        16'h68A8 : rd_rsp_data <= 32'h00000001;
        16'h6A20 : rd_rsp_data <= 32'h01000208;
        16'h6A24 : rd_rsp_data <= 32'h00000400;
        16'h6A28 : rd_rsp_data <= 32'h0100021A;
        16'h6A2C : rd_rsp_data <= 32'h00000400;
        16'h6A30 : rd_rsp_data <= 32'h0100021A;
        16'h6A34 : rd_rsp_data <= 32'h00000400;
        16'h6A38 : rd_rsp_data <= 32'h0100021A;
        16'h6A3C : rd_rsp_data <= 32'h00000C00;
        16'h6A40 : rd_rsp_data <= 32'h47000001;
        16'h6A48 : rd_rsp_data <= 32'h4B000001;
        16'h6A50 : rd_rsp_data <= 32'h47000001;
        16'h6A58 : rd_rsp_data <= 32'h4B000001;
        16'h6A60 : rd_rsp_data <= 32'h01000208;
        16'h6A64 : rd_rsp_data <= 32'h00000400;
        16'h6A68 : rd_rsp_data <= 32'h0100021A;
        16'h6A6C : rd_rsp_data <= 32'h00000400;
        16'h6B00 : rd_rsp_data <= 32'h01000208;
        16'h6B04 : rd_rsp_data <= 32'h00000400;
        16'h6B08 : rd_rsp_data <= 32'h0100020A;
        16'h6B0C : rd_rsp_data <= 32'h00000400;
        16'h6B10 : rd_rsp_data <= 32'h0100020A;
        16'h6B14 : rd_rsp_data <= 32'h00000400;
        16'h6C00 : rd_rsp_data <= 32'h00000003;
        16'h6C04 : rd_rsp_data <= 32'h50500101;
        16'h6C08 : rd_rsp_data <= 32'h84008300;
        16'h6C0C : rd_rsp_data <= 32'h01F10001;
        16'h6C10 : rd_rsp_data <= 32'h00000060;
        16'h6C14 : rd_rsp_data <= 32'h00000062;
        16'h6C1C : rd_rsp_data <= 32'h00000008;
        16'h6C2C : rd_rsp_data <= 32'h00F00000;
        16'h6C30 : rd_rsp_data <= 32'h0000FFF0;
        16'h6C34 : rd_rsp_data <= 32'h0001FFF1;
        16'h6C44 : rd_rsp_data <= 32'h0000000B;
        16'h6C54 : rd_rsp_data <= 32'h00F00000;
        16'h6C58 : rd_rsp_data <= 32'h0000FFF0;
        16'h6C5C : rd_rsp_data <= 32'h0001FFF1;
        16'h6C6C : rd_rsp_data <= 32'h0000000B;
        16'h6C80 : rd_rsp_data <= 32'h0000FFFF;
        16'h6C88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6C8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6C90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6C94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6C98 : rd_rsp_data <= 32'h00000001;
        16'h6C9C : rd_rsp_data <= 32'h0000FFFF;
        16'h6CA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6CA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6CA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6CAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6CB4 : rd_rsp_data <= 32'h00F00000;
        16'h6CB8 : rd_rsp_data <= 32'h0000FFF0;
        16'h6CBC : rd_rsp_data <= 32'h0001FFF1;
        16'h6CCC : rd_rsp_data <= 32'h00000008;
        16'h6CDC : rd_rsp_data <= 32'h00F00000;
        16'h6CE0 : rd_rsp_data <= 32'h0000FFF0;
        16'h6CE4 : rd_rsp_data <= 32'h0001FFF1;
        16'h6CF4 : rd_rsp_data <= 32'h00000008;
        16'h6D04 : rd_rsp_data <= 32'h00F00000;
        16'h6D08 : rd_rsp_data <= 32'h0000FFF0;
        16'h6D0C : rd_rsp_data <= 32'h0001FFF1;
        16'h6D1C : rd_rsp_data <= 32'h00000008;
        16'h6D2C : rd_rsp_data <= 32'h00F00000;
        16'h6D30 : rd_rsp_data <= 32'h0000FFF0;
        16'h6D34 : rd_rsp_data <= 32'h0001FFF1;
        16'h6D44 : rd_rsp_data <= 32'h00000008;
        16'h6D54 : rd_rsp_data <= 32'h00F00000;
        16'h6D58 : rd_rsp_data <= 32'h0000FFF0;
        16'h6D5C : rd_rsp_data <= 32'h0001FFF1;
        16'h6D6C : rd_rsp_data <= 32'h00000008;
        16'h6D7C : rd_rsp_data <= 32'h00F00000;
        16'h6D80 : rd_rsp_data <= 32'h0000FFF0;
        16'h6D84 : rd_rsp_data <= 32'h0001FFF1;
        16'h6D94 : rd_rsp_data <= 32'h00000008;
        16'h6DA4 : rd_rsp_data <= 32'h00F00000;
        16'h6DA8 : rd_rsp_data <= 32'h0000FFF0;
        16'h6DAC : rd_rsp_data <= 32'h0001FFF1;
        16'h6DBC : rd_rsp_data <= 32'h00000008;
        16'h6F30 : rd_rsp_data <= 32'h00000001;
        16'h6F40 : rd_rsp_data <= 32'h01101FF0;
        16'h6F44 : rd_rsp_data <= 32'h01200000;
        16'h6F48 : rd_rsp_data <= 32'h19001FE0;
        16'h6F4C : rd_rsp_data <= 32'h07000000;
        16'h6F50 : rd_rsp_data <= 32'hBDD683F9;
        16'h6F54 : rd_rsp_data <= 32'h0000000E;
        16'h6F58 : rd_rsp_data <= 32'hD5A1215F;
        16'h6F5C : rd_rsp_data <= 32'h0000000B;
        16'h6F60 : rd_rsp_data <= 32'h00000520;
        16'h6F70 : rd_rsp_data <= 32'hF73897F0;
        16'h6F74 : rd_rsp_data <= 32'h00000005;
        16'h6F80 : rd_rsp_data <= 32'h000000A4;
        16'h6F90 : rd_rsp_data <= 32'h19CFDB88;
        16'h6FA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6FA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6FAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6FB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h6FB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h7004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h7008 : rd_rsp_data <= 32'h800000F8;
        16'h7010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h7014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h7030 : rd_rsp_data <= 32'h000700B0;
        16'h7034 : rd_rsp_data <= 32'h000700B0;
        16'h7080 : rd_rsp_data <= 32'h01000208;
        16'h7084 : rd_rsp_data <= 32'h00000400;
        16'h7088 : rd_rsp_data <= 32'h0100030A;
        16'h708C : rd_rsp_data <= 32'h00000408;
        16'h7090 : rd_rsp_data <= 32'h00004000;
        16'h7094 : rd_rsp_data <= 32'h00011FFF;
        16'h7098 : rd_rsp_data <= 32'h00000060;
        16'h7100 : rd_rsp_data <= 32'h0810C008;
        16'h7110 : rd_rsp_data <= 32'hFB000001;
        16'h715C : rd_rsp_data <= 32'h00000001;
        16'h7160 : rd_rsp_data <= 32'h00000001;
        16'h7180 : rd_rsp_data <= 32'h01000208;
        16'h7184 : rd_rsp_data <= 32'h00000400;
        16'h7188 : rd_rsp_data <= 32'h0100021A;
        16'h718C : rd_rsp_data <= 32'h00000400;
        16'h7250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h7254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h725C : rd_rsp_data <= 32'h00000004;
        16'h7260 : rd_rsp_data <= 32'hAD7FFFFF;
        16'h7264 : rd_rsp_data <= 32'h00000004;
        16'h7268 : rd_rsp_data <= 32'h03082404;
        16'h7270 : rd_rsp_data <= 32'h00010000;
        16'h7278 : rd_rsp_data <= 32'h00000001;
        16'h7300 : rd_rsp_data <= 32'h00000023;
        16'h7400 : rd_rsp_data <= 32'h00000001;
        16'h7428 : rd_rsp_data <= 32'h000F0000;
        16'h7430 : rd_rsp_data <= 32'h41422484;
        16'h7434 : rd_rsp_data <= 32'h12416968;
        16'h7438 : rd_rsp_data <= 32'h41921888;
        16'h743C : rd_rsp_data <= 32'h12416918;
        16'h7444 : rd_rsp_data <= 32'h000000B0;
        16'h7450 : rd_rsp_data <= 32'h00060352;
        16'h7454 : rd_rsp_data <= 32'h0000020A;
        16'h7458 : rd_rsp_data <= 32'h0004A311;
        16'h745C : rd_rsp_data <= 32'h0000020A;
        16'h7460 : rd_rsp_data <= 32'h00048249;
        16'h7464 : rd_rsp_data <= 32'h00000209;
        16'h7468 : rd_rsp_data <= 32'h01C49249;
        16'h746C : rd_rsp_data <= 32'h00000209;
        16'h7470 : rd_rsp_data <= 32'h4C022D2A;
        16'h7474 : rd_rsp_data <= 32'h9BC24A21;
        16'h7478 : rd_rsp_data <= 32'h08308647;
        16'h747C : rd_rsp_data <= 32'h834241E1;
        16'h7480 : rd_rsp_data <= 32'h00049249;
        16'h7484 : rd_rsp_data <= 32'h00001209;
        16'h7488 : rd_rsp_data <= 32'h0F1009A5;
        16'h748C : rd_rsp_data <= 32'h6C0DC58F;
        16'h7490 : rd_rsp_data <= 32'h000010EF;
        16'h7498 : rd_rsp_data <= 32'h41921888;
        16'h749C : rd_rsp_data <= 32'h12416918;
        16'h74A0 : rd_rsp_data <= 32'h00000100;
        16'h74A4 : rd_rsp_data <= 32'h0000003F;
        16'h7500 : rd_rsp_data <= 32'h01010208;
        16'h7504 : rd_rsp_data <= 32'h00000400;
        16'h7510 : rd_rsp_data <= 32'h4101861F;
        16'h7514 : rd_rsp_data <= 32'h00001408;
        16'h7518 : rd_rsp_data <= 32'h0100021B;
        16'h751C : rd_rsp_data <= 32'h00000400;
        16'h7528 : rd_rsp_data <= 32'h0100021B;
        16'h752C : rd_rsp_data <= 32'h00000C00;
        16'h7530 : rd_rsp_data <= 32'h01000208;
        16'h7534 : rd_rsp_data <= 32'h00000400;
        16'h7538 : rd_rsp_data <= 32'h0100020A;
        16'h753C : rd_rsp_data <= 32'h00000400;
        16'h7540 : rd_rsp_data <= 32'h0100020A;
        16'h7544 : rd_rsp_data <= 32'h00000400;
        16'h7800 : rd_rsp_data <= 32'h00044400;
        16'h7804 : rd_rsp_data <= 32'h19321932;
        16'h7808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h780C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h7814 : rd_rsp_data <= 32'h000400BE;
        16'h7818 : rd_rsp_data <= 32'h000400BE;
        16'h782C : rd_rsp_data <= 32'h00000B63;
        16'h7854 : rd_rsp_data <= 32'h00842108;
        16'h7860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h7864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h7900 : rd_rsp_data <= 32'h0011C000;
        16'h7904 : rd_rsp_data <= 32'hFFFFC000;
        16'h7908 : rd_rsp_data <= 32'h01010210;
        16'h790C : rd_rsp_data <= 32'h00000400;
        16'h7910 : rd_rsp_data <= 32'h01010210;
        16'h7914 : rd_rsp_data <= 32'h00000400;
        16'h7918 : rd_rsp_data <= 32'h01010210;
        16'h791C : rd_rsp_data <= 32'h00000400;
        16'h7928 : rd_rsp_data <= 32'h01010210;
        16'h792C : rd_rsp_data <= 32'h00000400;
        16'h7930 : rd_rsp_data <= 32'h01010210;
        16'h7934 : rd_rsp_data <= 32'h00000400;
        16'h7938 : rd_rsp_data <= 32'h01010210;
        16'h793C : rd_rsp_data <= 32'h00000400;
        16'h7940 : rd_rsp_data <= 32'h00120000;
        16'h7944 : rd_rsp_data <= 32'hFFFFC000;
        16'h7948 : rd_rsp_data <= 32'h01010210;
        16'h794C : rd_rsp_data <= 32'h00000400;
        16'h7950 : rd_rsp_data <= 32'h01010210;
        16'h7954 : rd_rsp_data <= 32'h00020400;
        16'h7958 : rd_rsp_data <= 32'h01010210;
        16'h795C : rd_rsp_data <= 32'h00020400;
        16'h7968 : rd_rsp_data <= 32'h01010210;
        16'h796C : rd_rsp_data <= 32'h00000400;
        16'h7970 : rd_rsp_data <= 32'h01010210;
        16'h7974 : rd_rsp_data <= 32'h00000400;
        16'h7978 : rd_rsp_data <= 32'h01010210;
        16'h797C : rd_rsp_data <= 32'h00000400;
        16'h7988 : rd_rsp_data <= 32'h01010210;
        16'h798C : rd_rsp_data <= 32'h00000400;
        16'h7990 : rd_rsp_data <= 32'h01010210;
        16'h7994 : rd_rsp_data <= 32'h00000400;
        16'h7998 : rd_rsp_data <= 32'h01010210;
        16'h799C : rd_rsp_data <= 32'h00000400;
        16'h79A8 : rd_rsp_data <= 32'h01010210;
        16'h79AC : rd_rsp_data <= 32'h00000400;
        16'h79B0 : rd_rsp_data <= 32'h01010210;
        16'h79B4 : rd_rsp_data <= 32'h00000400;
        16'h79B8 : rd_rsp_data <= 32'h01010210;
        16'h79BC : rd_rsp_data <= 32'h00000400;
        16'h79C8 : rd_rsp_data <= 32'h01010210;
        16'h79CC : rd_rsp_data <= 32'h00000400;
        16'h79D0 : rd_rsp_data <= 32'h01010210;
        16'h79D4 : rd_rsp_data <= 32'h00000400;
        16'h79D8 : rd_rsp_data <= 32'h01010210;
        16'h79DC : rd_rsp_data <= 32'h00000400;
        16'h79E8 : rd_rsp_data <= 32'h01010210;
        16'h79EC : rd_rsp_data <= 32'h00000400;
        16'h79F0 : rd_rsp_data <= 32'h01010210;
        16'h79F4 : rd_rsp_data <= 32'h00000400;
        16'h79F8 : rd_rsp_data <= 32'h01010210;
        16'h79FC : rd_rsp_data <= 32'h00000400;
        16'h7A00 : rd_rsp_data <= 32'h00124000;
        16'h7A04 : rd_rsp_data <= 32'hFFFFF000;
        16'h7A08 : rd_rsp_data <= 32'h01010210;
        16'h7A0C : rd_rsp_data <= 32'h00000400;
        16'h7A10 : rd_rsp_data <= 32'h01000210;
        16'h7A14 : rd_rsp_data <= 32'h02000400;
        16'h7A18 : rd_rsp_data <= 32'h01000210;
        16'h7A1C : rd_rsp_data <= 32'h02000400;
        16'h7A28 : rd_rsp_data <= 32'h01010210;
        16'h7A2C : rd_rsp_data <= 32'h00000400;
        16'h7A30 : rd_rsp_data <= 32'h01010210;
        16'h7A34 : rd_rsp_data <= 32'h00000400;
        16'h7A38 : rd_rsp_data <= 32'h01010210;
        16'h7A3C : rd_rsp_data <= 32'h00000400;
        16'h7A48 : rd_rsp_data <= 32'h01010210;
        16'h7A4C : rd_rsp_data <= 32'h00000400;
        16'h7A50 : rd_rsp_data <= 32'h01010210;
        16'h7A54 : rd_rsp_data <= 32'h00000400;
        16'h7A58 : rd_rsp_data <= 32'h01010210;
        16'h7A5C : rd_rsp_data <= 32'h00000400;
        16'h7A68 : rd_rsp_data <= 32'h01010210;
        16'h7A6C : rd_rsp_data <= 32'h00000400;
        16'h7A70 : rd_rsp_data <= 32'h01010210;
        16'h7A74 : rd_rsp_data <= 32'h00000400;
        16'h7A78 : rd_rsp_data <= 32'h01010210;
        16'h7A7C : rd_rsp_data <= 32'h00000400;
        16'h7A80 : rd_rsp_data <= 32'h00125000;
        16'h7A84 : rd_rsp_data <= 32'hFFFFFFE0;
        16'h7A88 : rd_rsp_data <= 32'h01010210;
        16'h7A8C : rd_rsp_data <= 32'h00000400;
        16'h7A90 : rd_rsp_data <= 32'h01010210;
        16'h7A94 : rd_rsp_data <= 32'h00000400;
        16'h7A98 : rd_rsp_data <= 32'h01010210;
        16'h7A9C : rd_rsp_data <= 32'h00000400;
        16'h7AA8 : rd_rsp_data <= 32'h01000200;
        16'h7AAC : rd_rsp_data <= 32'h00000400;
        16'h7AC0 : rd_rsp_data <= 32'h00125020;
        16'h7AC4 : rd_rsp_data <= 32'hFFFFFFE0;
        16'h7AC8 : rd_rsp_data <= 32'h01010210;
        16'h7ACC : rd_rsp_data <= 32'h00000400;
        16'h7AD0 : rd_rsp_data <= 32'h01010210;
        16'h7AD4 : rd_rsp_data <= 32'h00000400;
        16'h7AD8 : rd_rsp_data <= 32'h01010210;
        16'h7ADC : rd_rsp_data <= 32'h00000400;
        16'h7AE0 : rd_rsp_data <= 32'h01000208;
        16'h7AE4 : rd_rsp_data <= 32'h00000400;
        16'h7AE8 : rd_rsp_data <= 32'h81000608;
        16'h7AEC : rd_rsp_data <= 32'h00001500;
        16'h7AF8 : rd_rsp_data <= 32'h01010210;
        16'h7AFC : rd_rsp_data <= 32'h00000400;
        16'h7B00 : rd_rsp_data <= 32'h01010210;
        16'h7B04 : rd_rsp_data <= 32'h00000400;
        16'h7B08 : rd_rsp_data <= 32'h01010210;
        16'h7B0C : rd_rsp_data <= 32'h00000400;
        16'h7B18 : rd_rsp_data <= 32'h01010210;
        16'h7B1C : rd_rsp_data <= 32'h00000400;
        16'h7B20 : rd_rsp_data <= 32'h01010210;
        16'h7B24 : rd_rsp_data <= 32'h00000400;
        16'h7B28 : rd_rsp_data <= 32'h01010210;
        16'h7B2C : rd_rsp_data <= 32'h00000400;
        16'h7B38 : rd_rsp_data <= 32'h01010210;
        16'h7B3C : rd_rsp_data <= 32'h00000400;
        16'h7B40 : rd_rsp_data <= 32'h01010210;
        16'h7B44 : rd_rsp_data <= 32'h00000400;
        16'h7B48 : rd_rsp_data <= 32'h01010210;
        16'h7B4C : rd_rsp_data <= 32'h00000400;
        16'h7B58 : rd_rsp_data <= 32'h01010210;
        16'h7B5C : rd_rsp_data <= 32'h00000400;
        16'h7B60 : rd_rsp_data <= 32'h01010210;
        16'h7B64 : rd_rsp_data <= 32'h00000400;
        16'h7B68 : rd_rsp_data <= 32'h01010210;
        16'h7B6C : rd_rsp_data <= 32'h00000400;
        16'h7B70 : rd_rsp_data <= 32'h00005105;
        16'h7B88 : rd_rsp_data <= 32'h01000208;
        16'h7B8C : rd_rsp_data <= 32'h00000400;
        16'h7B90 : rd_rsp_data <= 32'h0100021A;
        16'h7B94 : rd_rsp_data <= 32'h00000400;
        16'h8000 : rd_rsp_data <= 32'h00421D18;
        16'h8004 : rd_rsp_data <= 32'h002D0C0C;
        16'h8008 : rd_rsp_data <= 32'h003A1010;
        16'h800C : rd_rsp_data <= 32'h0025080C;
        16'h8010 : rd_rsp_data <= 32'h00351818;
        16'h8014 : rd_rsp_data <= 32'h00361818;
        16'h8018 : rd_rsp_data <= 32'h00182929;
        16'h801C : rd_rsp_data <= 32'h00351010;
        16'h8080 : rd_rsp_data <= 32'h10C68000;
        16'h8084 : rd_rsp_data <= 32'hF0F87843;
        16'h8088 : rd_rsp_data <= 32'hFC212480;
        16'h808C : rd_rsp_data <= 32'h005AC001;
        16'h8090 : rd_rsp_data <= 32'h4F9E1000;
        16'h8094 : rd_rsp_data <= 32'h00063C21;
        16'h8098 : rd_rsp_data <= 32'h4EE00000;
        16'h809C : rd_rsp_data <= 32'h0A025B81;
        16'h80A0 : rd_rsp_data <= 32'h9FF054FE;
        16'h80A4 : rd_rsp_data <= 32'h54210F76;
        16'h80A8 : rd_rsp_data <= 32'h98C011DF;
        16'h80AC : rd_rsp_data <= 32'hA8000000;
        16'h80B0 : rd_rsp_data <= 32'h045E4904;
        16'h80B4 : rd_rsp_data <= 32'h061C003B;
        16'h80B8 : rd_rsp_data <= 32'h8820EE1F;
        16'h80BC : rd_rsp_data <= 32'h58155D63;
        16'h80C8 : rd_rsp_data <= 32'h30000000;
        16'h80D4 : rd_rsp_data <= 32'h01041041;
        16'h80D8 : rd_rsp_data <= 32'h08208080;
        16'h80DC : rd_rsp_data <= 32'h1E560820;
        16'h80E0 : rd_rsp_data <= 32'h8062788B;
        16'h80E4 : rd_rsp_data <= 32'h745A6E72;
        16'h80E8 : rd_rsp_data <= 32'h80635C5C;
        16'h80EC : rd_rsp_data <= 32'h80808080;
        16'h80F0 : rd_rsp_data <= 32'h80808080;
        16'h80F4 : rd_rsp_data <= 32'h015AB343;
        16'h80F8 : rd_rsp_data <= 32'h01020FFF;
        16'h80FC : rd_rsp_data <= 32'h01020FFF;
        16'h8100 : rd_rsp_data <= 32'h01020FFF;
        16'h8108 : rd_rsp_data <= 32'h001D537F;
        16'h810C : rd_rsp_data <= 32'h00FFFFFF;
        16'h8110 : rd_rsp_data <= 32'h00FFFFFF;
        16'h8114 : rd_rsp_data <= 32'h00FFFFFF;
        16'h8128 : rd_rsp_data <= 32'h03800000;
        16'h812C : rd_rsp_data <= 32'h060D19EE;
        16'h813C : rd_rsp_data <= 32'h023200E5;
        16'h8140 : rd_rsp_data <= 32'h0006087E;
        16'h8148 : rd_rsp_data <= 32'h80100010;
        16'h814C : rd_rsp_data <= 32'h99999999;
        16'h8150 : rd_rsp_data <= 32'h210842F0;
        16'h8154 : rd_rsp_data <= 32'h210842F0;
        16'h8158 : rd_rsp_data <= 32'h210842B0;
        16'h815C : rd_rsp_data <= 32'h210842B0;
        16'h8160 : rd_rsp_data <= 32'h21084190;
        16'h8164 : rd_rsp_data <= 32'h210842B0;
        16'h8168 : rd_rsp_data <= 32'h21084270;
        16'h816C : rd_rsp_data <= 32'h21084210;
        16'h8170 : rd_rsp_data <= 32'h21084210;
        16'h8174 : rd_rsp_data <= 32'h21084210;
        16'h8178 : rd_rsp_data <= 32'h00084210;
        16'h817C : rd_rsp_data <= 32'h00077054;
        16'h8180 : rd_rsp_data <= 32'h08400000;
        16'h8198 : rd_rsp_data <= 32'h808CF60A;
        16'h819C : rd_rsp_data <= 32'h00000014;
        16'h81A0 : rd_rsp_data <= 32'h00019400;
        16'h81AC : rd_rsp_data <= 32'h03260244;
        16'h81B0 : rd_rsp_data <= 32'h12481000;
        16'h81B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h81B8 : rd_rsp_data <= 32'h05700036;
        16'h81BC : rd_rsp_data <= 32'h0154C222;
        16'h81C4 : rd_rsp_data <= 32'h000003F4;
        16'h81C8 : rd_rsp_data <= 32'h78000000;
        16'h81D8 : rd_rsp_data <= 32'h07400000;
        16'h81DC : rd_rsp_data <= 32'h02180080;
        16'h81E0 : rd_rsp_data <= 32'h00142000;
        16'h81E8 : rd_rsp_data <= 32'h40000000;
        16'h8200 : rd_rsp_data <= 32'h00322114;
        16'h8204 : rd_rsp_data <= 32'h00181810;
        16'h8208 : rd_rsp_data <= 32'h003E1C10;
        16'h820C : rd_rsp_data <= 32'h001C1818;
        16'h8210 : rd_rsp_data <= 32'h00101C18;
        16'h8214 : rd_rsp_data <= 32'h00281910;
        16'h8218 : rd_rsp_data <= 32'h00251414;
        16'h821C : rd_rsp_data <= 32'h00291008;
        16'h8280 : rd_rsp_data <= 32'h10C68000;
        16'h8284 : rd_rsp_data <= 32'hF0783801;
        16'h8288 : rd_rsp_data <= 32'hFC212480;
        16'h828C : rd_rsp_data <= 32'h005DC001;
        16'h8290 : rd_rsp_data <= 32'h4E9E1000;
        16'h8294 : rd_rsp_data <= 32'h00063C21;
        16'h8298 : rd_rsp_data <= 32'h5DE00000;
        16'h829C : rd_rsp_data <= 32'h0A025B81;
        16'h82A0 : rd_rsp_data <= 32'h9FF056FE;
        16'h82A4 : rd_rsp_data <= 32'hAC210F9E;
        16'h82A8 : rd_rsp_data <= 32'h98C011DF;
        16'h82AC : rd_rsp_data <= 32'hA8000000;
        16'h82B0 : rd_rsp_data <= 32'h045E4904;
        16'h82B4 : rd_rsp_data <= 32'h061C003B;
        16'h82B8 : rd_rsp_data <= 32'h8820EE1F;
        16'h82BC : rd_rsp_data <= 32'h58155D63;
        16'h82C8 : rd_rsp_data <= 32'h30000000;
        16'h82D4 : rd_rsp_data <= 32'h01041041;
        16'h82D8 : rd_rsp_data <= 32'h08208080;
        16'h82DC : rd_rsp_data <= 32'h1E560820;
        16'h82E0 : rd_rsp_data <= 32'h80624C8B;
        16'h82E4 : rd_rsp_data <= 32'h6E685F5C;
        16'h82E8 : rd_rsp_data <= 32'h80706966;
        16'h82EC : rd_rsp_data <= 32'h80808080;
        16'h82F0 : rd_rsp_data <= 32'h80808080;
        16'h82F4 : rd_rsp_data <= 32'h0162D2A1;
        16'h82F8 : rd_rsp_data <= 32'h01020FFF;
        16'h82FC : rd_rsp_data <= 32'h01020FFF;
        16'h8300 : rd_rsp_data <= 32'h01020FFF;
        16'h8308 : rd_rsp_data <= 32'h001C1363;
        16'h830C : rd_rsp_data <= 32'h00FFFFFF;
        16'h8310 : rd_rsp_data <= 32'h00FFFFFF;
        16'h8314 : rd_rsp_data <= 32'h00FFFFFF;
        16'h8320 : rd_rsp_data <= 32'h00006000;
        16'h8328 : rd_rsp_data <= 32'h03800000;
        16'h832C : rd_rsp_data <= 32'h064C1D7C;
        16'h833C : rd_rsp_data <= 32'h024204DC;
        16'h8340 : rd_rsp_data <= 32'h0006087E;
        16'h8348 : rd_rsp_data <= 32'h80100010;
        16'h834C : rd_rsp_data <= 32'h99999999;
        16'h8350 : rd_rsp_data <= 32'h21084210;
        16'h8354 : rd_rsp_data <= 32'h210842B0;
        16'h8358 : rd_rsp_data <= 32'h21084250;
        16'h835C : rd_rsp_data <= 32'h21084310;
        16'h8360 : rd_rsp_data <= 32'h21084210;
        16'h8364 : rd_rsp_data <= 32'h21084330;
        16'h8368 : rd_rsp_data <= 32'h21084270;
        16'h836C : rd_rsp_data <= 32'h21084230;
        16'h8370 : rd_rsp_data <= 32'h21084210;
        16'h8374 : rd_rsp_data <= 32'h21084210;
        16'h8378 : rd_rsp_data <= 32'h00084210;
        16'h837C : rd_rsp_data <= 32'h00077054;
        16'h8380 : rd_rsp_data <= 32'h08400000;
        16'h8398 : rd_rsp_data <= 32'h808CF60A;
        16'h839C : rd_rsp_data <= 32'h00000015;
        16'h83A0 : rd_rsp_data <= 32'h00019400;
        16'h83AC : rd_rsp_data <= 32'h03260244;
        16'h83B0 : rd_rsp_data <= 32'h12481000;
        16'h83B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h83B8 : rd_rsp_data <= 32'h05700036;
        16'h83BC : rd_rsp_data <= 32'h0154C222;
        16'h83C4 : rd_rsp_data <= 32'h000007A2;
        16'h83C8 : rd_rsp_data <= 32'h78900000;
        16'h83D8 : rd_rsp_data <= 32'h07400000;
        16'h83DC : rd_rsp_data <= 32'h02180080;
        16'h83E0 : rd_rsp_data <= 32'h00152000;
        16'h83E8 : rd_rsp_data <= 32'h40000000;
        16'h8400 : rd_rsp_data <= 32'h00421D18;
        16'h8404 : rd_rsp_data <= 32'h002D0C0C;
        16'h8408 : rd_rsp_data <= 32'h003A1010;
        16'h840C : rd_rsp_data <= 32'h0025080C;
        16'h8410 : rd_rsp_data <= 32'h00351818;
        16'h8414 : rd_rsp_data <= 32'h00361818;
        16'h8418 : rd_rsp_data <= 32'h00182929;
        16'h841C : rd_rsp_data <= 32'h00351010;
        16'h8480 : rd_rsp_data <= 32'h10C68000;
        16'h8484 : rd_rsp_data <= 32'hF0F87843;
        16'h8488 : rd_rsp_data <= 32'hFC212480;
        16'h848C : rd_rsp_data <= 32'h005AC001;
        16'h8490 : rd_rsp_data <= 32'h4F9E1000;
        16'h8494 : rd_rsp_data <= 32'h00063C21;
        16'h8498 : rd_rsp_data <= 32'h4EE00000;
        16'h849C : rd_rsp_data <= 32'h0A025B81;
        16'h84A0 : rd_rsp_data <= 32'h9FF054FE;
        16'h84A4 : rd_rsp_data <= 32'h54210F76;
        16'h84A8 : rd_rsp_data <= 32'h98C011DF;
        16'h84AC : rd_rsp_data <= 32'hA8000000;
        16'h84B0 : rd_rsp_data <= 32'h045E4904;
        16'h84B4 : rd_rsp_data <= 32'h061C003B;
        16'h84B8 : rd_rsp_data <= 32'h8820EE1F;
        16'h84BC : rd_rsp_data <= 32'h58155D63;
        16'h84C8 : rd_rsp_data <= 32'h30000000;
        16'h84D4 : rd_rsp_data <= 32'h01041041;
        16'h84D8 : rd_rsp_data <= 32'h08208080;
        16'h84DC : rd_rsp_data <= 32'h1E560820;
        16'h84E0 : rd_rsp_data <= 32'h8062788B;
        16'h84E4 : rd_rsp_data <= 32'h745A6E72;
        16'h84E8 : rd_rsp_data <= 32'h80635C5C;
        16'h84EC : rd_rsp_data <= 32'h80808080;
        16'h84F0 : rd_rsp_data <= 32'h80808080;
        16'h84F4 : rd_rsp_data <= 32'h015AB343;
        16'h84F8 : rd_rsp_data <= 32'h01020FFF;
        16'h84FC : rd_rsp_data <= 32'h01020FFF;
        16'h8500 : rd_rsp_data <= 32'h01020FFF;
        16'h8508 : rd_rsp_data <= 32'h001D537F;
        16'h850C : rd_rsp_data <= 32'h00FFFFFF;
        16'h8510 : rd_rsp_data <= 32'h00FFFFFF;
        16'h8514 : rd_rsp_data <= 32'h00FFFFFF;
        16'h8528 : rd_rsp_data <= 32'h03800000;
        16'h852C : rd_rsp_data <= 32'h060D19EE;
        16'h853C : rd_rsp_data <= 32'h023200E5;
        16'h8540 : rd_rsp_data <= 32'h0006087E;
        16'h8548 : rd_rsp_data <= 32'h80100010;
        16'h854C : rd_rsp_data <= 32'h99999999;
        16'h8550 : rd_rsp_data <= 32'h210842F0;
        16'h8554 : rd_rsp_data <= 32'h210842F0;
        16'h8558 : rd_rsp_data <= 32'h210842B0;
        16'h855C : rd_rsp_data <= 32'h210842B0;
        16'h8560 : rd_rsp_data <= 32'h21084190;
        16'h8564 : rd_rsp_data <= 32'h210842B0;
        16'h8568 : rd_rsp_data <= 32'h21084270;
        16'h856C : rd_rsp_data <= 32'h21084210;
        16'h8570 : rd_rsp_data <= 32'h21084210;
        16'h8574 : rd_rsp_data <= 32'h21084210;
        16'h8578 : rd_rsp_data <= 32'h00084210;
        16'h857C : rd_rsp_data <= 32'h00077054;
        16'h8580 : rd_rsp_data <= 32'h08400000;
        16'h8598 : rd_rsp_data <= 32'h808CF60A;
        16'h859C : rd_rsp_data <= 32'h00000014;
        16'h85A0 : rd_rsp_data <= 32'h00019400;
        16'h85AC : rd_rsp_data <= 32'h03260244;
        16'h85B0 : rd_rsp_data <= 32'h12481000;
        16'h85B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h85B8 : rd_rsp_data <= 32'h05700036;
        16'h85BC : rd_rsp_data <= 32'h0154C222;
        16'h85C4 : rd_rsp_data <= 32'h000003F4;
        16'h85C8 : rd_rsp_data <= 32'h78000000;
        16'h85D8 : rd_rsp_data <= 32'h07400000;
        16'h85DC : rd_rsp_data <= 32'h02180080;
        16'h85E0 : rd_rsp_data <= 32'h00142000;
        16'h85E8 : rd_rsp_data <= 32'h40000000;
        16'h8600 : rd_rsp_data <= 32'h2001FC0B;
        16'h8604 : rd_rsp_data <= 32'h00000005;
        16'h8608 : rd_rsp_data <= 32'h009C0000;
        16'h860C : rd_rsp_data <= 32'h00800092;
        16'h8610 : rd_rsp_data <= 32'h00000100;
        16'h8614 : rd_rsp_data <= 32'h00000080;
        16'h8618 : rd_rsp_data <= 32'h057E4804;
        16'h861C : rd_rsp_data <= 32'h0000003B;
        16'h8620 : rd_rsp_data <= 32'h8020F207;
        16'h8624 : rd_rsp_data <= 32'h40155D63;
        16'h8628 : rd_rsp_data <= 32'h00000075;
        16'h862C : rd_rsp_data <= 32'h3FFE0000;
        16'h8630 : rd_rsp_data <= 32'h0000020F;
        16'h863C : rd_rsp_data <= 32'h60E7D545;
        16'h8640 : rd_rsp_data <= 32'h0005C478;
        16'h8648 : rd_rsp_data <= 32'h0E400010;
        16'h8658 : rd_rsp_data <= 32'h0F000000;
        16'h8660 : rd_rsp_data <= 32'h808F8887;
        16'h8664 : rd_rsp_data <= 32'h9B918F7C;
        16'h8668 : rd_rsp_data <= 32'h8B89918B;
        16'h866C : rd_rsp_data <= 32'hFF94899C;
        16'h8670 : rd_rsp_data <= 32'h80808080;
        16'h8674 : rd_rsp_data <= 32'h98902001;
        16'h8680 : rd_rsp_data <= 32'h00E20000;
        16'h8688 : rd_rsp_data <= 32'h00000006;
        16'h868C : rd_rsp_data <= 32'h0001CA00;
        16'h8690 : rd_rsp_data <= 32'h01660444;
        16'h8694 : rd_rsp_data <= 32'hE00DCE0C;
        16'h869C : rd_rsp_data <= 32'h08400000;
        16'h86B4 : rd_rsp_data <= 32'h07500000;
        16'h86B8 : rd_rsp_data <= 32'h82A885DC;
        16'h86BC : rd_rsp_data <= 32'h027816A0;
        16'h86C0 : rd_rsp_data <= 32'h02C2061D;
        16'h86C4 : rd_rsp_data <= 32'h0154C222;
        16'h86CC : rd_rsp_data <= 32'h01440000;
        16'h86D0 : rd_rsp_data <= 32'hFFFF0000;
        16'h86D4 : rd_rsp_data <= 32'h20000000;
        16'h86FC : rd_rsp_data <= 32'h00062000;
        16'h8700 : rd_rsp_data <= 32'h2001FC0B;
        16'h8704 : rd_rsp_data <= 32'h00000005;
        16'h8708 : rd_rsp_data <= 32'h009E0000;
        16'h870C : rd_rsp_data <= 32'h00800094;
        16'h8710 : rd_rsp_data <= 32'h00000100;
        16'h8714 : rd_rsp_data <= 32'h00000080;
        16'h8718 : rd_rsp_data <= 32'h057E4804;
        16'h871C : rd_rsp_data <= 32'h0000003B;
        16'h8720 : rd_rsp_data <= 32'h8020E207;
        16'h8724 : rd_rsp_data <= 32'h40155D63;
        16'h8728 : rd_rsp_data <= 32'h00000075;
        16'h872C : rd_rsp_data <= 32'h3FFE0000;
        16'h8730 : rd_rsp_data <= 32'h0000020F;
        16'h873C : rd_rsp_data <= 32'h60E7D545;
        16'h8740 : rd_rsp_data <= 32'h0005C478;
        16'h8748 : rd_rsp_data <= 32'h0E400010;
        16'h8758 : rd_rsp_data <= 32'h0F000000;
        16'h8760 : rd_rsp_data <= 32'h808D7887;
        16'h8764 : rd_rsp_data <= 32'h7C89888C;
        16'h8768 : rd_rsp_data <= 32'h78808D7C;
        16'h876C : rd_rsp_data <= 32'hFF90857C;
        16'h8770 : rd_rsp_data <= 32'h80808080;
        16'h8774 : rd_rsp_data <= 32'h89852001;
        16'h8780 : rd_rsp_data <= 32'h00E20000;
        16'h8788 : rd_rsp_data <= 32'h00000006;
        16'h878C : rd_rsp_data <= 32'h0001CA00;
        16'h8790 : rd_rsp_data <= 32'h01660444;
        16'h8794 : rd_rsp_data <= 32'hE00DCE0C;
        16'h879C : rd_rsp_data <= 32'h08400000;
        16'h87B4 : rd_rsp_data <= 32'h07500000;
        16'h87B8 : rd_rsp_data <= 32'h82A885DC;
        16'h87BC : rd_rsp_data <= 32'h027816A0;
        16'h87C0 : rd_rsp_data <= 32'h02C2061D;
        16'h87C4 : rd_rsp_data <= 32'h0154C222;
        16'h87CC : rd_rsp_data <= 32'h01440000;
        16'h87D0 : rd_rsp_data <= 32'hFFFF0000;
        16'h87D4 : rd_rsp_data <= 32'h20000000;
        16'h87E8 : rd_rsp_data <= 32'h000005EC;
        16'h87FC : rd_rsp_data <= 32'h00062000;
        16'h8800 : rd_rsp_data <= 32'h2001FC0B;
        16'h8804 : rd_rsp_data <= 32'h00000005;
        16'h8808 : rd_rsp_data <= 32'h009C0000;
        16'h880C : rd_rsp_data <= 32'h00800092;
        16'h8810 : rd_rsp_data <= 32'h00000100;
        16'h8814 : rd_rsp_data <= 32'h00000080;
        16'h8818 : rd_rsp_data <= 32'h057E4804;
        16'h881C : rd_rsp_data <= 32'h0000003B;
        16'h8820 : rd_rsp_data <= 32'h8020F207;
        16'h8824 : rd_rsp_data <= 32'h40155D63;
        16'h8828 : rd_rsp_data <= 32'h00000075;
        16'h882C : rd_rsp_data <= 32'h3FFE0000;
        16'h8830 : rd_rsp_data <= 32'h0000020F;
        16'h883C : rd_rsp_data <= 32'h60E7D545;
        16'h8840 : rd_rsp_data <= 32'h0005C478;
        16'h8848 : rd_rsp_data <= 32'h0E400010;
        16'h8858 : rd_rsp_data <= 32'h0F000000;
        16'h8860 : rd_rsp_data <= 32'h808F8887;
        16'h8864 : rd_rsp_data <= 32'h9B918F7C;
        16'h8868 : rd_rsp_data <= 32'h8B89918B;
        16'h886C : rd_rsp_data <= 32'hFF94899C;
        16'h8870 : rd_rsp_data <= 32'h80808080;
        16'h8874 : rd_rsp_data <= 32'h98902001;
        16'h8880 : rd_rsp_data <= 32'h00E20000;
        16'h8888 : rd_rsp_data <= 32'h00000006;
        16'h888C : rd_rsp_data <= 32'h0001CA00;
        16'h8890 : rd_rsp_data <= 32'h01660444;
        16'h8894 : rd_rsp_data <= 32'hE00DCE0C;
        16'h889C : rd_rsp_data <= 32'h08400000;
        16'h88B4 : rd_rsp_data <= 32'h07500000;
        16'h88B8 : rd_rsp_data <= 32'h82A885DC;
        16'h88BC : rd_rsp_data <= 32'h027816A0;
        16'h88C0 : rd_rsp_data <= 32'h02C2061D;
        16'h88C4 : rd_rsp_data <= 32'h0154C222;
        16'h88CC : rd_rsp_data <= 32'h01440000;
        16'h88D0 : rd_rsp_data <= 32'hFFFF0000;
        16'h88D4 : rd_rsp_data <= 32'h20000000;
        16'h88FC : rd_rsp_data <= 32'h00062000;
        16'h8900 : rd_rsp_data <= 32'h2001FC0B;
        16'h8904 : rd_rsp_data <= 32'h00000005;
        16'h8908 : rd_rsp_data <= 32'h009E0000;
        16'h890C : rd_rsp_data <= 32'h00800094;
        16'h8910 : rd_rsp_data <= 32'h00000100;
        16'h8914 : rd_rsp_data <= 32'h00000080;
        16'h8918 : rd_rsp_data <= 32'h057E4804;
        16'h891C : rd_rsp_data <= 32'h0000003B;
        16'h8920 : rd_rsp_data <= 32'h8020E207;
        16'h8924 : rd_rsp_data <= 32'h40155D63;
        16'h8928 : rd_rsp_data <= 32'h00000075;
        16'h892C : rd_rsp_data <= 32'h3FFE0000;
        16'h8930 : rd_rsp_data <= 32'h0000020F;
        16'h893C : rd_rsp_data <= 32'h60E7D545;
        16'h8940 : rd_rsp_data <= 32'h0005C478;
        16'h8948 : rd_rsp_data <= 32'h0E400010;
        16'h8958 : rd_rsp_data <= 32'h0F000000;
        16'h8960 : rd_rsp_data <= 32'h808D7887;
        16'h8964 : rd_rsp_data <= 32'h7C89888C;
        16'h8968 : rd_rsp_data <= 32'h78808D7C;
        16'h896C : rd_rsp_data <= 32'hFF90857C;
        16'h8970 : rd_rsp_data <= 32'h80808080;
        16'h8974 : rd_rsp_data <= 32'h89852001;
        16'h8980 : rd_rsp_data <= 32'h00E20000;
        16'h8988 : rd_rsp_data <= 32'h00000006;
        16'h898C : rd_rsp_data <= 32'h0001CA00;
        16'h8990 : rd_rsp_data <= 32'h01660444;
        16'h8994 : rd_rsp_data <= 32'hE00DCE0C;
        16'h899C : rd_rsp_data <= 32'h08400000;
        16'h89B4 : rd_rsp_data <= 32'h07500000;
        16'h89B8 : rd_rsp_data <= 32'h82A885DC;
        16'h89BC : rd_rsp_data <= 32'h027816A0;
        16'h89C0 : rd_rsp_data <= 32'h02C2061D;
        16'h89C4 : rd_rsp_data <= 32'h0154C222;
        16'h89CC : rd_rsp_data <= 32'h01440000;
        16'h89D0 : rd_rsp_data <= 32'hFFFF0000;
        16'h89D4 : rd_rsp_data <= 32'h20000000;
        16'h89E8 : rd_rsp_data <= 32'h000005EC;
        16'h89FC : rd_rsp_data <= 32'h00062000;
        16'h8A00 : rd_rsp_data <= 32'h2001F590;
        16'h8A04 : rd_rsp_data <= 32'h00000005;
        16'h8A08 : rd_rsp_data <= 32'h007E0000;
        16'h8A0C : rd_rsp_data <= 32'h00800080;
        16'h8A10 : rd_rsp_data <= 32'h00000100;
        16'h8A18 : rd_rsp_data <= 32'h057E4804;
        16'h8A1C : rd_rsp_data <= 32'h0000003B;
        16'h8A20 : rd_rsp_data <= 32'h8020E607;
        16'h8A24 : rd_rsp_data <= 32'h40155D63;
        16'h8A28 : rd_rsp_data <= 32'h00000075;
        16'h8A2C : rd_rsp_data <= 32'h3FFE0000;
        16'h8A30 : rd_rsp_data <= 32'h0000020F;
        16'h8A3C : rd_rsp_data <= 32'h60E7D545;
        16'h8A40 : rd_rsp_data <= 32'h0005C478;
        16'h8A48 : rd_rsp_data <= 32'h0E400010;
        16'h8A58 : rd_rsp_data <= 32'h0F000000;
        16'h8A60 : rd_rsp_data <= 32'h80928F68;
        16'h8A64 : rd_rsp_data <= 32'h87909094;
        16'h8A68 : rd_rsp_data <= 32'h89878185;
        16'h8A6C : rd_rsp_data <= 32'hFF909089;
        16'h8A70 : rd_rsp_data <= 32'h80808080;
        16'h8A74 : rd_rsp_data <= 32'h7C802001;
        16'h8A80 : rd_rsp_data <= 32'h00E20000;
        16'h8A88 : rd_rsp_data <= 32'h00000006;
        16'h8A8C : rd_rsp_data <= 32'h0001CA00;
        16'h8A90 : rd_rsp_data <= 32'h01660444;
        16'h8A94 : rd_rsp_data <= 32'hE00DCE0C;
        16'h8A9C : rd_rsp_data <= 32'h08400000;
        16'h8AB4 : rd_rsp_data <= 32'h07500000;
        16'h8AB8 : rd_rsp_data <= 32'h82A885DC;
        16'h8ABC : rd_rsp_data <= 32'h027816A0;
        16'h8AC0 : rd_rsp_data <= 32'h02C2061D;
        16'h8AC4 : rd_rsp_data <= 32'h0154C222;
        16'h8ACC : rd_rsp_data <= 32'h01440000;
        16'h8AD0 : rd_rsp_data <= 32'hFFFF0000;
        16'h8AD4 : rd_rsp_data <= 32'h20000000;
        16'h8AE8 : rd_rsp_data <= 32'h0000037C;
        16'h8AFC : rd_rsp_data <= 32'h00062000;
        16'h8B00 : rd_rsp_data <= 32'h2001FC0B;
        16'h8B04 : rd_rsp_data <= 32'h00000005;
        16'h8B08 : rd_rsp_data <= 32'h009C0000;
        16'h8B0C : rd_rsp_data <= 32'h00800092;
        16'h8B10 : rd_rsp_data <= 32'h00000100;
        16'h8B14 : rd_rsp_data <= 32'h00000080;
        16'h8B18 : rd_rsp_data <= 32'h057E4804;
        16'h8B1C : rd_rsp_data <= 32'h0000003B;
        16'h8B20 : rd_rsp_data <= 32'h8020F207;
        16'h8B24 : rd_rsp_data <= 32'h40155D63;
        16'h8B28 : rd_rsp_data <= 32'h00000075;
        16'h8B2C : rd_rsp_data <= 32'h3FFE0000;
        16'h8B30 : rd_rsp_data <= 32'h0000020F;
        16'h8B3C : rd_rsp_data <= 32'h60E7D545;
        16'h8B40 : rd_rsp_data <= 32'h0005C478;
        16'h8B48 : rd_rsp_data <= 32'h0E400010;
        16'h8B58 : rd_rsp_data <= 32'h0F000000;
        16'h8B60 : rd_rsp_data <= 32'h808F8887;
        16'h8B64 : rd_rsp_data <= 32'h9B918F7C;
        16'h8B68 : rd_rsp_data <= 32'h8B89918B;
        16'h8B6C : rd_rsp_data <= 32'hFF94899C;
        16'h8B70 : rd_rsp_data <= 32'h80808080;
        16'h8B74 : rd_rsp_data <= 32'h98902001;
        16'h8B80 : rd_rsp_data <= 32'h00E20000;
        16'h8B88 : rd_rsp_data <= 32'h00000006;
        16'h8B8C : rd_rsp_data <= 32'h0001CA00;
        16'h8B90 : rd_rsp_data <= 32'h01660444;
        16'h8B94 : rd_rsp_data <= 32'hE00DCE0C;
        16'h8B9C : rd_rsp_data <= 32'h08400000;
        16'h8BB4 : rd_rsp_data <= 32'h07500000;
        16'h8BB8 : rd_rsp_data <= 32'h82A885DC;
        16'h8BBC : rd_rsp_data <= 32'h027816A0;
        16'h8BC0 : rd_rsp_data <= 32'h02C2061D;
        16'h8BC4 : rd_rsp_data <= 32'h0154C222;
        16'h8BCC : rd_rsp_data <= 32'h01440000;
        16'h8BD0 : rd_rsp_data <= 32'hFFFF0000;
        16'h8BD4 : rd_rsp_data <= 32'h20000000;
        16'h8BFC : rd_rsp_data <= 32'h00062000;
        16'h8C00 : rd_rsp_data <= 32'h00000003;
        16'h8C08 : rd_rsp_data <= 32'h0640E9A0;
        16'h8C10 : rd_rsp_data <= 32'h3BFBEFBD;
        16'h8C14 : rd_rsp_data <= 32'h0000003E;
        16'h8C18 : rd_rsp_data <= 32'h00000001;
        16'h8C80 : rd_rsp_data <= 32'h00000001;
        16'h8C84 : rd_rsp_data <= 32'h000C3C3C;
        16'h8C8C : rd_rsp_data <= 32'h00000001;
        16'h8C90 : rd_rsp_data <= 32'h17171D1D;
        16'h8C9C : rd_rsp_data <= 32'h190F1622;
        16'h8CA0 : rd_rsp_data <= 32'h052AAAD1;
        16'h8D00 : rd_rsp_data <= 32'h00001503;
        16'h8D04 : rd_rsp_data <= 32'h00FF0F0F;
        16'h8D08 : rd_rsp_data <= 32'h00082315;
        16'h8D80 : rd_rsp_data <= 32'h000C3C3C;
        16'h8D8C : rd_rsp_data <= 32'h00000001;
        16'h8D90 : rd_rsp_data <= 32'h50000000;
        16'h8D94 : rd_rsp_data <= 32'h60C02000;
        16'h8DA0 : rd_rsp_data <= 32'h08600080;
        16'h8DA4 : rd_rsp_data <= 32'h08600080;
        16'h8DB0 : rd_rsp_data <= 32'hFCF1DEF0;
        16'h8DB4 : rd_rsp_data <= 32'hFF7DCE7C;
        16'h8DB8 : rd_rsp_data <= 32'hE7F7B000;
        16'h8DBC : rd_rsp_data <= 32'h110F1622;
        16'h8DC0 : rd_rsp_data <= 32'h0B44A555;
        16'h8DC4 : rd_rsp_data <= 32'h007AC72B;
        16'h8DC8 : rd_rsp_data <= 32'h00000D3B;
        16'h8E00 : rd_rsp_data <= 32'h2001F470;
        16'h8E04 : rd_rsp_data <= 32'h00000005;
        16'h8E08 : rd_rsp_data <= 32'h00820000;
        16'h8E0C : rd_rsp_data <= 32'h00800080;
        16'h8E10 : rd_rsp_data <= 32'h00000100;
        16'h8E18 : rd_rsp_data <= 32'h057E4804;
        16'h8E1C : rd_rsp_data <= 32'h0000003B;
        16'h8E20 : rd_rsp_data <= 32'h8020F207;
        16'h8E24 : rd_rsp_data <= 32'h40155D63;
        16'h8E28 : rd_rsp_data <= 32'h00000075;
        16'h8E2C : rd_rsp_data <= 32'h3FFE0000;
        16'h8E30 : rd_rsp_data <= 32'h0000020F;
        16'h8E3C : rd_rsp_data <= 32'h60E7D545;
        16'h8E40 : rd_rsp_data <= 32'h0005C478;
        16'h8E48 : rd_rsp_data <= 32'h0E400010;
        16'h8E58 : rd_rsp_data <= 32'h0F000000;
        16'h8E60 : rd_rsp_data <= 32'h80939478;
        16'h8E64 : rd_rsp_data <= 32'h7C9C918F;
        16'h8E68 : rd_rsp_data <= 32'h9885857E;
        16'h8E6C : rd_rsp_data <= 32'hFF94919F;
        16'h8E70 : rd_rsp_data <= 32'h80808080;
        16'h8E74 : rd_rsp_data <= 32'h93982001;
        16'h8E80 : rd_rsp_data <= 32'h00E20000;
        16'h8E8C : rd_rsp_data <= 32'h0001CA00;
        16'h8E90 : rd_rsp_data <= 32'h01660444;
        16'h8E94 : rd_rsp_data <= 32'hE00DCE0C;
        16'h8E9C : rd_rsp_data <= 32'h08400000;
        16'h8EB4 : rd_rsp_data <= 32'h07500000;
        16'h8EB8 : rd_rsp_data <= 32'h82A885DC;
        16'h8EBC : rd_rsp_data <= 32'h027816A0;
        16'h8EC0 : rd_rsp_data <= 32'h02C2061D;
        16'h8EC4 : rd_rsp_data <= 32'h0154C222;
        16'h8ECC : rd_rsp_data <= 32'h01440000;
        16'h8ED0 : rd_rsp_data <= 32'hFFFF0000;
        16'h8ED4 : rd_rsp_data <= 32'h20000000;
        16'h8EFC : rd_rsp_data <= 32'h00002000;
        16'h8F00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8F9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h8FFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h900C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h901C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h902C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h903C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h904C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h905C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h906C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h907C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h908C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h909C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h90FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h910C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h911C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h912C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h913C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h914C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h915C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h916C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h917C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h918C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h919C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h91FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9200 : rd_rsp_data <= 32'h000C0C08;
        16'h9204 : rd_rsp_data <= 32'h0029100C;
        16'h9208 : rd_rsp_data <= 32'h00100C08;
        16'h920C : rd_rsp_data <= 32'h00180C04;
        16'h9210 : rd_rsp_data <= 32'h0021140C;
        16'h9214 : rd_rsp_data <= 32'h001C100C;
        16'h9218 : rd_rsp_data <= 32'h00081410;
        16'h921C : rd_rsp_data <= 32'h00181910;
        16'h9280 : rd_rsp_data <= 32'h10C68000;
        16'h9284 : rd_rsp_data <= 32'hF0F87843;
        16'h9288 : rd_rsp_data <= 32'hFC212480;
        16'h928C : rd_rsp_data <= 32'h0057C001;
        16'h9290 : rd_rsp_data <= 32'h4F9E1000;
        16'h9294 : rd_rsp_data <= 32'h00063C21;
        16'h9298 : rd_rsp_data <= 32'h4FE00000;
        16'h929C : rd_rsp_data <= 32'h0A025B81;
        16'h92A0 : rd_rsp_data <= 32'h9FF0573E;
        16'h92A4 : rd_rsp_data <= 32'h54210FBF;
        16'h92A8 : rd_rsp_data <= 32'h98C011DF;
        16'h92AC : rd_rsp_data <= 32'hA8000000;
        16'h92B0 : rd_rsp_data <= 32'h045E4904;
        16'h92B4 : rd_rsp_data <= 32'h061C003B;
        16'h92B8 : rd_rsp_data <= 32'h8820E21F;
        16'h92BC : rd_rsp_data <= 32'h58155D63;
        16'h92C8 : rd_rsp_data <= 32'h30000000;
        16'h92D4 : rd_rsp_data <= 32'h01041041;
        16'h92D8 : rd_rsp_data <= 32'h08208080;
        16'h92DC : rd_rsp_data <= 32'h1E560820;
        16'h92E0 : rd_rsp_data <= 32'h80627078;
        16'h92E4 : rd_rsp_data <= 32'h504A645D;
        16'h92E8 : rd_rsp_data <= 32'h806C6B68;
        16'h92EC : rd_rsp_data <= 32'h80808080;
        16'h92F0 : rd_rsp_data <= 32'h80808080;
        16'h92F4 : rd_rsp_data <= 32'h0142C3FD;
        16'h92F8 : rd_rsp_data <= 32'h01020FFF;
        16'h92FC : rd_rsp_data <= 32'h01020FFF;
        16'h9300 : rd_rsp_data <= 32'h01020FFF;
        16'h9308 : rd_rsp_data <= 32'h002093C1;
        16'h930C : rd_rsp_data <= 32'h00FFFFFF;
        16'h9310 : rd_rsp_data <= 32'h00FFFFFF;
        16'h9314 : rd_rsp_data <= 32'h00FFFFFF;
        16'h9320 : rd_rsp_data <= 32'h0001D000;
        16'h9328 : rd_rsp_data <= 32'h03800000;
        16'h932C : rd_rsp_data <= 32'h07458BBC;
        16'h933C : rd_rsp_data <= 32'h023600E3;
        16'h9340 : rd_rsp_data <= 32'h0006087E;
        16'h9348 : rd_rsp_data <= 32'h80100010;
        16'h934C : rd_rsp_data <= 32'h99999999;
        16'h9350 : rd_rsp_data <= 32'h21084210;
        16'h9354 : rd_rsp_data <= 32'h21084210;
        16'h9358 : rd_rsp_data <= 32'h210841F0;
        16'h935C : rd_rsp_data <= 32'h21084210;
        16'h9360 : rd_rsp_data <= 32'h21084270;
        16'h9364 : rd_rsp_data <= 32'h21084270;
        16'h9368 : rd_rsp_data <= 32'h21084250;
        16'h936C : rd_rsp_data <= 32'h21084270;
        16'h9370 : rd_rsp_data <= 32'h21084210;
        16'h9374 : rd_rsp_data <= 32'h21084210;
        16'h9378 : rd_rsp_data <= 32'h00084210;
        16'h937C : rd_rsp_data <= 32'h00077054;
        16'h9380 : rd_rsp_data <= 32'h08400000;
        16'h9398 : rd_rsp_data <= 32'h808CF60A;
        16'h939C : rd_rsp_data <= 32'h00000016;
        16'h93A0 : rd_rsp_data <= 32'h00019400;
        16'h93AC : rd_rsp_data <= 32'h03260244;
        16'h93B0 : rd_rsp_data <= 32'h12481000;
        16'h93B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h93B8 : rd_rsp_data <= 32'h05700036;
        16'h93BC : rd_rsp_data <= 32'h0154C222;
        16'h93C4 : rd_rsp_data <= 32'h00000754;
        16'h93C8 : rd_rsp_data <= 32'h78000000;
        16'h93D8 : rd_rsp_data <= 32'h07400000;
        16'h93DC : rd_rsp_data <= 32'h02180080;
        16'h93E0 : rd_rsp_data <= 32'h00162000;
        16'h93E8 : rd_rsp_data <= 32'h40000000;
        16'h9400 : rd_rsp_data <= 32'h00421D18;
        16'h9404 : rd_rsp_data <= 32'h002D0C0C;
        16'h9408 : rd_rsp_data <= 32'h003A1010;
        16'h940C : rd_rsp_data <= 32'h0025080C;
        16'h9410 : rd_rsp_data <= 32'h00351818;
        16'h9414 : rd_rsp_data <= 32'h00361818;
        16'h9418 : rd_rsp_data <= 32'h00182929;
        16'h941C : rd_rsp_data <= 32'h00351010;
        16'h9480 : rd_rsp_data <= 32'h11C680A0;
        16'h9484 : rd_rsp_data <= 32'hF0F87843;
        16'h9488 : rd_rsp_data <= 32'hFC212480;
        16'h948C : rd_rsp_data <= 32'h005AC001;
        16'h9490 : rd_rsp_data <= 32'h4FDE1800;
        16'h9494 : rd_rsp_data <= 32'h00063C63;
        16'h9498 : rd_rsp_data <= 32'h4EE00000;
        16'h949C : rd_rsp_data <= 32'h0A03DB81;
        16'h94A0 : rd_rsp_data <= 32'h9FF077FE;
        16'h94A4 : rd_rsp_data <= 32'hD4210FFF;
        16'h94A8 : rd_rsp_data <= 32'hD8C011DF;
        16'h94AC : rd_rsp_data <= 32'hA8000000;
        16'h94B0 : rd_rsp_data <= 32'h045E6904;
        16'h94B4 : rd_rsp_data <= 32'h061D023B;
        16'h94B8 : rd_rsp_data <= 32'h8820EE1F;
        16'h94BC : rd_rsp_data <= 32'h5817FDE7;
        16'h94C8 : rd_rsp_data <= 32'h38000000;
        16'h94D4 : rd_rsp_data <= 32'h01041041;
        16'h94D8 : rd_rsp_data <= 32'h08209090;
        16'h94DC : rd_rsp_data <= 32'h3E7E0820;
        16'h94E0 : rd_rsp_data <= 32'h80E2F88B;
        16'h94E4 : rd_rsp_data <= 32'hF4DAEEF2;
        16'h94E8 : rd_rsp_data <= 32'h80E3DCDC;
        16'h94EC : rd_rsp_data <= 32'h80808080;
        16'h94F0 : rd_rsp_data <= 32'h80808080;
        16'h94F4 : rd_rsp_data <= 32'h015ABFFF;
        16'h94F8 : rd_rsp_data <= 32'h01020FFF;
        16'h94FC : rd_rsp_data <= 32'h01020FFF;
        16'h9500 : rd_rsp_data <= 32'h01020FFF;
        16'h9508 : rd_rsp_data <= 32'h00FFFFFF;
        16'h950C : rd_rsp_data <= 32'h00FFFFFF;
        16'h9510 : rd_rsp_data <= 32'h00FFFFFF;
        16'h9514 : rd_rsp_data <= 32'h00FFFFFF;
        16'h9528 : rd_rsp_data <= 32'h03800000;
        16'h952C : rd_rsp_data <= 32'h06FFDFEE;
        16'h953C : rd_rsp_data <= 32'h023200E5;
        16'h9540 : rd_rsp_data <= 32'h0006087E;
        16'h9548 : rd_rsp_data <= 32'h80100010;
        16'h954C : rd_rsp_data <= 32'h99999999;
        16'h9550 : rd_rsp_data <= 32'h210842F0;
        16'h9554 : rd_rsp_data <= 32'h210842F0;
        16'h9558 : rd_rsp_data <= 32'h210842B0;
        16'h955C : rd_rsp_data <= 32'h210842B0;
        16'h9560 : rd_rsp_data <= 32'h21084390;
        16'h9564 : rd_rsp_data <= 32'h210842B0;
        16'h9568 : rd_rsp_data <= 32'h21084270;
        16'h956C : rd_rsp_data <= 32'h21084210;
        16'h9570 : rd_rsp_data <= 32'h21084210;
        16'h9574 : rd_rsp_data <= 32'h21084210;
        16'h9578 : rd_rsp_data <= 32'h00084210;
        16'h957C : rd_rsp_data <= 32'h00077254;
        16'h9580 : rd_rsp_data <= 32'h08400000;
        16'h9598 : rd_rsp_data <= 32'h808CF60A;
        16'h959C : rd_rsp_data <= 32'h00000414;
        16'h95A0 : rd_rsp_data <= 32'h00019400;
        16'h95AC : rd_rsp_data <= 32'h03260244;
        16'h95B0 : rd_rsp_data <= 32'h12481000;
        16'h95B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h95B8 : rd_rsp_data <= 32'h05700036;
        16'h95BC : rd_rsp_data <= 32'h0154C222;
        16'h95C4 : rd_rsp_data <= 32'h000007FE;
        16'h95C8 : rd_rsp_data <= 32'h78000000;
        16'h95D8 : rd_rsp_data <= 32'h07400000;
        16'h95DC : rd_rsp_data <= 32'h02180080;
        16'h95E0 : rd_rsp_data <= 32'h00142000;
        16'h95E8 : rd_rsp_data <= 32'h40000000;
        16'h9600 : rd_rsp_data <= 32'h000C0C08;
        16'h9604 : rd_rsp_data <= 32'h0029100C;
        16'h9608 : rd_rsp_data <= 32'h00100C08;
        16'h960C : rd_rsp_data <= 32'h00180C04;
        16'h9610 : rd_rsp_data <= 32'h0021140C;
        16'h9614 : rd_rsp_data <= 32'h001C100C;
        16'h9618 : rd_rsp_data <= 32'h00081410;
        16'h961C : rd_rsp_data <= 32'h00181910;
        16'h9680 : rd_rsp_data <= 32'h10C68000;
        16'h9684 : rd_rsp_data <= 32'hF0F87843;
        16'h9688 : rd_rsp_data <= 32'hFC212480;
        16'h968C : rd_rsp_data <= 32'h0057C001;
        16'h9690 : rd_rsp_data <= 32'h4F9E1000;
        16'h9694 : rd_rsp_data <= 32'h00063C21;
        16'h9698 : rd_rsp_data <= 32'h4FE00000;
        16'h969C : rd_rsp_data <= 32'h0A025B81;
        16'h96A0 : rd_rsp_data <= 32'h9FF0573E;
        16'h96A4 : rd_rsp_data <= 32'h54210FBF;
        16'h96A8 : rd_rsp_data <= 32'h98C011DF;
        16'h96AC : rd_rsp_data <= 32'hA8000000;
        16'h96B0 : rd_rsp_data <= 32'h045E4904;
        16'h96B4 : rd_rsp_data <= 32'h061C003B;
        16'h96B8 : rd_rsp_data <= 32'h8820E21F;
        16'h96BC : rd_rsp_data <= 32'h58155D63;
        16'h96C8 : rd_rsp_data <= 32'h30000000;
        16'h96D4 : rd_rsp_data <= 32'h01041041;
        16'h96D8 : rd_rsp_data <= 32'h08208080;
        16'h96DC : rd_rsp_data <= 32'h1E560820;
        16'h96E0 : rd_rsp_data <= 32'h80627078;
        16'h96E4 : rd_rsp_data <= 32'h504A645D;
        16'h96E8 : rd_rsp_data <= 32'h806C6B68;
        16'h96EC : rd_rsp_data <= 32'h80808080;
        16'h96F0 : rd_rsp_data <= 32'h80808080;
        16'h96F4 : rd_rsp_data <= 32'h0142C3FD;
        16'h96F8 : rd_rsp_data <= 32'h01020FFF;
        16'h96FC : rd_rsp_data <= 32'h01020FFF;
        16'h9700 : rd_rsp_data <= 32'h01020FFF;
        16'h9708 : rd_rsp_data <= 32'h002093C1;
        16'h970C : rd_rsp_data <= 32'h00FFFFFF;
        16'h9710 : rd_rsp_data <= 32'h00FFFFFF;
        16'h9714 : rd_rsp_data <= 32'h00FFFFFF;
        16'h9720 : rd_rsp_data <= 32'h0001D000;
        16'h9728 : rd_rsp_data <= 32'h03800000;
        16'h972C : rd_rsp_data <= 32'h07458BBC;
        16'h973C : rd_rsp_data <= 32'h023600E3;
        16'h9740 : rd_rsp_data <= 32'h0006087E;
        16'h9748 : rd_rsp_data <= 32'h80100010;
        16'h974C : rd_rsp_data <= 32'h99999999;
        16'h9750 : rd_rsp_data <= 32'h21084210;
        16'h9754 : rd_rsp_data <= 32'h21084210;
        16'h9758 : rd_rsp_data <= 32'h210841F0;
        16'h975C : rd_rsp_data <= 32'h21084210;
        16'h9760 : rd_rsp_data <= 32'h21084270;
        16'h9764 : rd_rsp_data <= 32'h21084270;
        16'h9768 : rd_rsp_data <= 32'h21084250;
        16'h976C : rd_rsp_data <= 32'h21084270;
        16'h9770 : rd_rsp_data <= 32'h21084210;
        16'h9774 : rd_rsp_data <= 32'h21084210;
        16'h9778 : rd_rsp_data <= 32'h00084210;
        16'h977C : rd_rsp_data <= 32'h00077054;
        16'h9780 : rd_rsp_data <= 32'h08400000;
        16'h9798 : rd_rsp_data <= 32'h808CF60A;
        16'h979C : rd_rsp_data <= 32'h00000016;
        16'h97A0 : rd_rsp_data <= 32'h00019400;
        16'h97AC : rd_rsp_data <= 32'h03260244;
        16'h97B0 : rd_rsp_data <= 32'h12481000;
        16'h97B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h97B8 : rd_rsp_data <= 32'h05700036;
        16'h97BC : rd_rsp_data <= 32'h0154C222;
        16'h97C4 : rd_rsp_data <= 32'h00000754;
        16'h97C8 : rd_rsp_data <= 32'h78000000;
        16'h97D8 : rd_rsp_data <= 32'h07400000;
        16'h97DC : rd_rsp_data <= 32'h02180080;
        16'h97E0 : rd_rsp_data <= 32'h00162000;
        16'h97E8 : rd_rsp_data <= 32'h40000000;
        16'h9800 : rd_rsp_data <= 32'h00421D18;
        16'h9804 : rd_rsp_data <= 32'h002D0C0C;
        16'h9808 : rd_rsp_data <= 32'h003A1010;
        16'h980C : rd_rsp_data <= 32'h0025080C;
        16'h9810 : rd_rsp_data <= 32'h00351818;
        16'h9814 : rd_rsp_data <= 32'h00361818;
        16'h9818 : rd_rsp_data <= 32'h00182929;
        16'h981C : rd_rsp_data <= 32'h00351010;
        16'h9880 : rd_rsp_data <= 32'h10C68000;
        16'h9884 : rd_rsp_data <= 32'hF0F87843;
        16'h9888 : rd_rsp_data <= 32'hFC212480;
        16'h988C : rd_rsp_data <= 32'h005AC001;
        16'h9890 : rd_rsp_data <= 32'h4F9E1000;
        16'h9894 : rd_rsp_data <= 32'h00063C21;
        16'h9898 : rd_rsp_data <= 32'h4EE00000;
        16'h989C : rd_rsp_data <= 32'h0A025B81;
        16'h98A0 : rd_rsp_data <= 32'h9FF054FE;
        16'h98A4 : rd_rsp_data <= 32'h54210F76;
        16'h98A8 : rd_rsp_data <= 32'h98C011DF;
        16'h98AC : rd_rsp_data <= 32'hA8000000;
        16'h98B0 : rd_rsp_data <= 32'h045E4904;
        16'h98B4 : rd_rsp_data <= 32'h061C003B;
        16'h98B8 : rd_rsp_data <= 32'h8820EE1F;
        16'h98BC : rd_rsp_data <= 32'h58155D63;
        16'h98C8 : rd_rsp_data <= 32'h30000000;
        16'h98D4 : rd_rsp_data <= 32'h01041041;
        16'h98D8 : rd_rsp_data <= 32'h08208080;
        16'h98DC : rd_rsp_data <= 32'h1E560820;
        16'h98E0 : rd_rsp_data <= 32'h8062788B;
        16'h98E4 : rd_rsp_data <= 32'h745A6E72;
        16'h98E8 : rd_rsp_data <= 32'h80635C5C;
        16'h98EC : rd_rsp_data <= 32'h80808080;
        16'h98F0 : rd_rsp_data <= 32'h80808080;
        16'h98F4 : rd_rsp_data <= 32'h015AB343;
        16'h98F8 : rd_rsp_data <= 32'h01020FFF;
        16'h98FC : rd_rsp_data <= 32'h01020FFF;
        16'h9900 : rd_rsp_data <= 32'h01020FFF;
        16'h9908 : rd_rsp_data <= 32'h001D537F;
        16'h990C : rd_rsp_data <= 32'h00FFFFFF;
        16'h9910 : rd_rsp_data <= 32'h00FFFFFF;
        16'h9914 : rd_rsp_data <= 32'h00FFFFFF;
        16'h9928 : rd_rsp_data <= 32'h03800000;
        16'h992C : rd_rsp_data <= 32'h060D19EE;
        16'h993C : rd_rsp_data <= 32'h023200E5;
        16'h9940 : rd_rsp_data <= 32'h0006087E;
        16'h9948 : rd_rsp_data <= 32'h80100010;
        16'h994C : rd_rsp_data <= 32'h99999999;
        16'h9950 : rd_rsp_data <= 32'h210842F0;
        16'h9954 : rd_rsp_data <= 32'h210842F0;
        16'h9958 : rd_rsp_data <= 32'h210842B0;
        16'h995C : rd_rsp_data <= 32'h210842B0;
        16'h9960 : rd_rsp_data <= 32'h21084190;
        16'h9964 : rd_rsp_data <= 32'h210842B0;
        16'h9968 : rd_rsp_data <= 32'h21084270;
        16'h996C : rd_rsp_data <= 32'h21084210;
        16'h9970 : rd_rsp_data <= 32'h21084210;
        16'h9974 : rd_rsp_data <= 32'h21084210;
        16'h9978 : rd_rsp_data <= 32'h00084210;
        16'h997C : rd_rsp_data <= 32'h00077054;
        16'h9980 : rd_rsp_data <= 32'h08400000;
        16'h9998 : rd_rsp_data <= 32'h808CF60A;
        16'h999C : rd_rsp_data <= 32'h00000014;
        16'h99A0 : rd_rsp_data <= 32'h00019400;
        16'h99AC : rd_rsp_data <= 32'h03260244;
        16'h99B0 : rd_rsp_data <= 32'h12481000;
        16'h99B4 : rd_rsp_data <= 32'h2D495C3E;
        16'h99B8 : rd_rsp_data <= 32'h05700036;
        16'h99BC : rd_rsp_data <= 32'h0154C222;
        16'h99C4 : rd_rsp_data <= 32'h000003F4;
        16'h99C8 : rd_rsp_data <= 32'h78000000;
        16'h99D8 : rd_rsp_data <= 32'h07400000;
        16'h99DC : rd_rsp_data <= 32'h02180080;
        16'h99E0 : rd_rsp_data <= 32'h00142000;
        16'h99E8 : rd_rsp_data <= 32'h40000000;
        16'h9A00 : rd_rsp_data <= 32'h001C1414;
        16'h9A04 : rd_rsp_data <= 32'h00311414;
        16'h9A08 : rd_rsp_data <= 32'h00081819;
        16'h9A0C : rd_rsp_data <= 32'h0024181C;
        16'h9A10 : rd_rsp_data <= 32'h00211D1D;
        16'h9A14 : rd_rsp_data <= 32'h00100C0C;
        16'h9A18 : rd_rsp_data <= 32'h001D181C;
        16'h9A1C : rd_rsp_data <= 32'h000C1418;
        16'h9A80 : rd_rsp_data <= 32'h10C68000;
        16'h9A84 : rd_rsp_data <= 32'hF0F87843;
        16'h9A88 : rd_rsp_data <= 32'hFC212480;
        16'h9A8C : rd_rsp_data <= 32'h0053C001;
        16'h9A90 : rd_rsp_data <= 32'h4F1E1000;
        16'h9A94 : rd_rsp_data <= 32'h00063C21;
        16'h9A98 : rd_rsp_data <= 32'h4FE00000;
        16'h9A9C : rd_rsp_data <= 32'h0A025B81;
        16'h9AA0 : rd_rsp_data <= 32'h9FF0577E;
        16'h9AA4 : rd_rsp_data <= 32'h1C210FBE;
        16'h9AA8 : rd_rsp_data <= 32'h98C011DF;
        16'h9AAC : rd_rsp_data <= 32'hA8000000;
        16'h9AB0 : rd_rsp_data <= 32'h045E4904;
        16'h9AB4 : rd_rsp_data <= 32'h061C003B;
        16'h9AB8 : rd_rsp_data <= 32'h8820E21F;
        16'h9ABC : rd_rsp_data <= 32'h58155D63;
        16'h9AC8 : rd_rsp_data <= 32'h30000000;
        16'h9AD4 : rd_rsp_data <= 32'h01041041;
        16'h9AD8 : rd_rsp_data <= 32'h08208080;
        16'h9ADC : rd_rsp_data <= 32'h1E560820;
        16'h9AE0 : rd_rsp_data <= 32'h806D4D93;
        16'h9AE4 : rd_rsp_data <= 32'h68646467;
        16'h9AE8 : rd_rsp_data <= 32'h80525A56;
        16'h9AEC : rd_rsp_data <= 32'h80808080;
        16'h9AF0 : rd_rsp_data <= 32'h80808080;
        16'h9AF4 : rd_rsp_data <= 32'h01429339;
        16'h9AF8 : rd_rsp_data <= 32'h01020FFF;
        16'h9AFC : rd_rsp_data <= 32'h01020FFF;
        16'h9B00 : rd_rsp_data <= 32'h01020FFF;
        16'h9B08 : rd_rsp_data <= 32'h001F13AB;
        16'h9B0C : rd_rsp_data <= 32'h00FFFFFF;
        16'h9B10 : rd_rsp_data <= 32'h00FFFFFF;
        16'h9B14 : rd_rsp_data <= 32'h00FFFFFF;
        16'h9B20 : rd_rsp_data <= 32'h0001A000;
        16'h9B28 : rd_rsp_data <= 32'h03800000;
        16'h9B2C : rd_rsp_data <= 32'h076889AF;
        16'h9B3C : rd_rsp_data <= 32'h023004E3;
        16'h9B40 : rd_rsp_data <= 32'h0006087E;
        16'h9B48 : rd_rsp_data <= 32'h80100010;
        16'h9B4C : rd_rsp_data <= 32'h99999999;
        16'h9B50 : rd_rsp_data <= 32'h21084290;
        16'h9B54 : rd_rsp_data <= 32'h210842D0;
        16'h9B58 : rd_rsp_data <= 32'h21084230;
        16'h9B5C : rd_rsp_data <= 32'h210841F0;
        16'h9B60 : rd_rsp_data <= 32'h21084270;
        16'h9B64 : rd_rsp_data <= 32'h21084250;
        16'h9B68 : rd_rsp_data <= 32'h21084250;
        16'h9B6C : rd_rsp_data <= 32'h21084250;
        16'h9B70 : rd_rsp_data <= 32'h21084210;
        16'h9B74 : rd_rsp_data <= 32'h21084210;
        16'h9B78 : rd_rsp_data <= 32'h00084210;
        16'h9B7C : rd_rsp_data <= 32'h00077054;
        16'h9B80 : rd_rsp_data <= 32'h08400000;
        16'h9B98 : rd_rsp_data <= 32'h808CF60A;
        16'h9B9C : rd_rsp_data <= 32'h00000016;
        16'h9BA0 : rd_rsp_data <= 32'h00019400;
        16'h9BAC : rd_rsp_data <= 32'h03260244;
        16'h9BB0 : rd_rsp_data <= 32'h12481000;
        16'h9BB4 : rd_rsp_data <= 32'h2D495C3E;
        16'h9BB8 : rd_rsp_data <= 32'h05700036;
        16'h9BBC : rd_rsp_data <= 32'h0154C222;
        16'h9BC4 : rd_rsp_data <= 32'h0000076E;
        16'h9BC8 : rd_rsp_data <= 32'h78000000;
        16'h9BD8 : rd_rsp_data <= 32'h07400000;
        16'h9BDC : rd_rsp_data <= 32'h02180080;
        16'h9BE0 : rd_rsp_data <= 32'h00162000;
        16'h9BE8 : rd_rsp_data <= 32'h40000000;
        16'h9C00 : rd_rsp_data <= 32'h00322114;
        16'h9C04 : rd_rsp_data <= 32'h00181810;
        16'h9C08 : rd_rsp_data <= 32'h003E1C10;
        16'h9C0C : rd_rsp_data <= 32'h001C1818;
        16'h9C10 : rd_rsp_data <= 32'h00101C18;
        16'h9C14 : rd_rsp_data <= 32'h00281910;
        16'h9C18 : rd_rsp_data <= 32'h00251414;
        16'h9C1C : rd_rsp_data <= 32'h00291008;
        16'h9C80 : rd_rsp_data <= 32'h10C68000;
        16'h9C84 : rd_rsp_data <= 32'hF0783801;
        16'h9C88 : rd_rsp_data <= 32'hFC212480;
        16'h9C8C : rd_rsp_data <= 32'h005DC001;
        16'h9C90 : rd_rsp_data <= 32'h4E9E1000;
        16'h9C94 : rd_rsp_data <= 32'h00063C21;
        16'h9C98 : rd_rsp_data <= 32'h5DE00000;
        16'h9C9C : rd_rsp_data <= 32'h0A025B81;
        16'h9CA0 : rd_rsp_data <= 32'h9FF056FE;
        16'h9CA4 : rd_rsp_data <= 32'hAC210F9E;
        16'h9CA8 : rd_rsp_data <= 32'h98C011DF;
        16'h9CAC : rd_rsp_data <= 32'hA8000000;
        16'h9CB0 : rd_rsp_data <= 32'h045E4904;
        16'h9CB4 : rd_rsp_data <= 32'h061C003B;
        16'h9CB8 : rd_rsp_data <= 32'h8820EE1F;
        16'h9CBC : rd_rsp_data <= 32'h58155D63;
        16'h9CC8 : rd_rsp_data <= 32'h30000000;
        16'h9CD4 : rd_rsp_data <= 32'h01041041;
        16'h9CD8 : rd_rsp_data <= 32'h08208080;
        16'h9CDC : rd_rsp_data <= 32'h1E560820;
        16'h9CE0 : rd_rsp_data <= 32'h80624C8B;
        16'h9CE4 : rd_rsp_data <= 32'h6E685F5C;
        16'h9CE8 : rd_rsp_data <= 32'h80706966;
        16'h9CEC : rd_rsp_data <= 32'h80808080;
        16'h9CF0 : rd_rsp_data <= 32'h80808080;
        16'h9CF4 : rd_rsp_data <= 32'h0162D2A1;
        16'h9CF8 : rd_rsp_data <= 32'h01020FFF;
        16'h9CFC : rd_rsp_data <= 32'h01020FFF;
        16'h9D00 : rd_rsp_data <= 32'h01020FFF;
        16'h9D08 : rd_rsp_data <= 32'h001C1363;
        16'h9D0C : rd_rsp_data <= 32'h00FFFFFF;
        16'h9D10 : rd_rsp_data <= 32'h00FFFFFF;
        16'h9D14 : rd_rsp_data <= 32'h00FFFFFF;
        16'h9D20 : rd_rsp_data <= 32'h00006000;
        16'h9D28 : rd_rsp_data <= 32'h03800000;
        16'h9D2C : rd_rsp_data <= 32'h064C1D7C;
        16'h9D3C : rd_rsp_data <= 32'h024204DC;
        16'h9D40 : rd_rsp_data <= 32'h0006087E;
        16'h9D48 : rd_rsp_data <= 32'h80100010;
        16'h9D4C : rd_rsp_data <= 32'h99999999;
        16'h9D50 : rd_rsp_data <= 32'h21084210;
        16'h9D54 : rd_rsp_data <= 32'h210842B0;
        16'h9D58 : rd_rsp_data <= 32'h21084250;
        16'h9D5C : rd_rsp_data <= 32'h21084310;
        16'h9D60 : rd_rsp_data <= 32'h21084210;
        16'h9D64 : rd_rsp_data <= 32'h21084330;
        16'h9D68 : rd_rsp_data <= 32'h21084270;
        16'h9D6C : rd_rsp_data <= 32'h21084230;
        16'h9D70 : rd_rsp_data <= 32'h21084210;
        16'h9D74 : rd_rsp_data <= 32'h21084210;
        16'h9D78 : rd_rsp_data <= 32'h00084210;
        16'h9D7C : rd_rsp_data <= 32'h00077054;
        16'h9D80 : rd_rsp_data <= 32'h08400000;
        16'h9D98 : rd_rsp_data <= 32'h808CF60A;
        16'h9D9C : rd_rsp_data <= 32'h00000015;
        16'h9DA0 : rd_rsp_data <= 32'h00019400;
        16'h9DAC : rd_rsp_data <= 32'h03260244;
        16'h9DB0 : rd_rsp_data <= 32'h12481000;
        16'h9DB4 : rd_rsp_data <= 32'h2D495C3E;
        16'h9DB8 : rd_rsp_data <= 32'h05700036;
        16'h9DBC : rd_rsp_data <= 32'h0154C222;
        16'h9DC4 : rd_rsp_data <= 32'h000007A2;
        16'h9DC8 : rd_rsp_data <= 32'h7F000000;
        16'h9DD8 : rd_rsp_data <= 32'h07400000;
        16'h9DDC : rd_rsp_data <= 32'h02180080;
        16'h9DE0 : rd_rsp_data <= 32'h00152000;
        16'h9DE8 : rd_rsp_data <= 32'h40000000;
        16'h9E00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9E9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9ECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9ED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9ED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9ED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9EFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h9F00 : rd_rsp_data <= 32'h0001860E;
        16'h9F04 : rd_rsp_data <= 32'h00015820;
        16'h9F0C : rd_rsp_data <= 32'h6C820008;
        16'h9F10 : rd_rsp_data <= 32'h00000402;
        16'h9F14 : rd_rsp_data <= 32'h3B000001;
        16'h9F18 : rd_rsp_data <= 32'hC1B20022;
        16'h9F1C : rd_rsp_data <= 32'h00410000;
        16'h9F20 : rd_rsp_data <= 32'h00000100;
        16'h9F24 : rd_rsp_data <= 32'h10003001;
        16'h9F28 : rd_rsp_data <= 32'h10100000;
        16'h9F2C : rd_rsp_data <= 32'h0010E2C0;
        16'h9F30 : rd_rsp_data <= 32'h1831BD44;
        16'h9F34 : rd_rsp_data <= 32'h0182B060;
        16'h9F38 : rd_rsp_data <= 32'hC0040534;
        16'h9F3C : rd_rsp_data <= 32'h602AD500;
        16'h9F40 : rd_rsp_data <= 32'hE0D50000;
        16'h9F48 : rd_rsp_data <= 32'h13004000;
        16'h9F4C : rd_rsp_data <= 32'h3C130E40;
        16'h9F50 : rd_rsp_data <= 32'h0145930E;
        16'h9F54 : rd_rsp_data <= 32'hFCD068AD;
        16'h9F58 : rd_rsp_data <= 32'h6C9B3062;
        16'h9F5C : rd_rsp_data <= 32'h00000001;
        16'h9F60 : rd_rsp_data <= 32'h1C104457;
        16'h9F64 : rd_rsp_data <= 32'h00006C82;
        16'h9F6C : rd_rsp_data <= 32'h04000000;
        16'h9F70 : rd_rsp_data <= 32'h00A8C754;
        16'h9F74 : rd_rsp_data <= 32'h0000C756;
        16'h9FA0 : rd_rsp_data <= 32'h00000908;
        16'h9FC4 : rd_rsp_data <= 32'h00000400;
        16'h9FC8 : rd_rsp_data <= 32'h00000001;
        16'h9FCC : rd_rsp_data <= 32'h000004E4;
        16'h9FD4 : rd_rsp_data <= 32'h00000001;
        16'h9FD8 : rd_rsp_data <= 32'h47200000;
        16'hA080 : rd_rsp_data <= 32'h08400000;
        16'hA098 : rd_rsp_data <= 32'h808CF60A;
        16'hA09C : rd_rsp_data <= 32'h00000415;
        16'hA0A0 : rd_rsp_data <= 32'h00019400;
        16'hA0AC : rd_rsp_data <= 32'h03260244;
        16'hA0B0 : rd_rsp_data <= 32'h12481000;
        16'hA0B4 : rd_rsp_data <= 32'h2D495C3E;
        16'hA0B8 : rd_rsp_data <= 32'h05700036;
        16'hA0BC : rd_rsp_data <= 32'h0154C222;
        16'hA0C4 : rd_rsp_data <= 32'h000007FE;
        16'hA0C8 : rd_rsp_data <= 32'h78000000;
        16'hA0D8 : rd_rsp_data <= 32'h07400000;
        16'hA0DC : rd_rsp_data <= 32'h02180080;
        16'hA0E0 : rd_rsp_data <= 32'h00152000;
        16'hA0E8 : rd_rsp_data <= 32'h40000000;
        16'hA100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA10C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA11C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA12C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA13C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA14C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA15C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA16C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA17C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA18C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA19C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA1FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA20C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA21C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA22C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA23C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA24C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA25C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA26C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA27C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA28C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA29C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA2FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA30C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA31C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA32C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA33C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA34C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA35C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA36C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA37C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA38C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA39C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA3FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA40C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA41C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA42C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA43C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA44C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA45C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA46C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA47C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA48C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA49C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA4FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA50C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA51C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA52C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA53C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA54C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA55C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA56C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA57C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA58C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA59C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA5FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA60C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA61C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA62C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA63C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA64C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA65C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA66C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA67C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA68C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA69C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA6FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA70C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA71C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA72C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA73C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA74C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA75C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA76C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA77C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA78C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA79C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA7FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA80C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA81C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA82C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA83C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA84C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA85C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA86C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA87C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA88C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA89C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA8FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA90C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA91C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA92C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA93C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA94C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA95C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA96C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA97C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA98C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA99C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hA9FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAA9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAAFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAB9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hABFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAC9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hACFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAD9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hADFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAE9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAEFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAF9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hAFFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB00C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB01C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB02C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB03C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB04C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB05C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB06C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB07C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB08C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB09C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB0FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB10C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB11C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB12C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB13C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB14C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB15C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB16C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB17C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB18C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB19C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB1FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB20C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB21C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB22C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB23C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB24C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB25C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB26C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB27C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB28C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB29C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB2FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB30C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB31C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB32C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB33C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB34C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB35C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB36C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB37C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB38C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB39C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB3FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB40C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB41C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB42C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB43C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB44C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB45C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB46C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB47C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB48C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB49C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB4FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB50C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB51C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB52C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB53C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB54C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB55C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB56C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB57C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB58C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB59C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB5FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB60C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB61C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB62C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB63C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB64C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB65C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB66C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB67C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB68C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB69C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB6FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB70C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB71C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB72C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB73C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB74C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB75C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB76C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB77C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB78C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB79C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB7FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB80C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB81C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB82C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB83C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB84C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB85C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB86C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB87C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB88C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB89C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB8FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB90C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB91C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB92C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB93C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB94C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB95C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB96C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB97C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB98C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB99C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hB9FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBA9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBAFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBB9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBBFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBC9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBCFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBD9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBDFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBE9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBEFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBF9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hBFFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC00C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC01C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC02C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC03C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC04C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC05C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC06C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC07C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC08C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC09C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC0FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC10C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC11C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC12C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC13C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC14C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC15C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC16C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC17C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC18C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC19C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC1FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC20C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC21C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC22C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC23C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC24C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC25C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC26C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC27C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC28C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC29C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC2FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC30C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC31C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC32C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC33C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC34C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC35C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC36C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC37C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC38C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC39C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC3FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC40C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC41C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC42C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC43C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC44C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC45C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC46C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC47C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC48C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC49C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC4FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC50C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC51C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC52C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC53C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC54C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC55C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC56C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC57C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC58C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC59C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC5FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC60C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC61C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC62C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC63C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC64C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC65C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC66C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC67C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC68C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC69C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC6FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC70C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC71C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC72C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC73C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC74C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC75C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC76C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC77C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC78C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC79C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC7FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC80C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC81C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC82C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC83C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC84C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC85C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC86C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC87C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC88C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC89C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC8FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC90C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC91C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC92C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC93C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC94C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC95C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC96C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC97C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC98C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC99C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hC9FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCA9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCAFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCB9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCBFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCC9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCCFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCD9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCDFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCE9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCEFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCF9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hCFFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD000 : rd_rsp_data <= 32'h01000208;
        16'hD004 : rd_rsp_data <= 32'h00000400;
        16'hD008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD00C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD010 : rd_rsp_data <= 32'h0100021A;
        16'hD014 : rd_rsp_data <= 32'h00000400;
        16'hD01C : rd_rsp_data <= 32'h00001800;
        16'hD028 : rd_rsp_data <= 32'h01040000;
        16'hD030 : rd_rsp_data <= 32'h00411421;
        16'hD038 : rd_rsp_data <= 32'h00010101;
        16'hD040 : rd_rsp_data <= 32'h0000AA55;
        16'hD044 : rd_rsp_data <= 32'h0000AA55;
        16'hD048 : rd_rsp_data <= 32'h0000AA55;
        16'hD050 : rd_rsp_data <= 32'h01010100;
        16'hD058 : rd_rsp_data <= 32'h80000000;
        16'hD05C : rd_rsp_data <= 32'h80000000;
        16'hD060 : rd_rsp_data <= 32'h80000000;
        16'hD100 : rd_rsp_data <= 32'h01000208;
        16'hD104 : rd_rsp_data <= 32'h00000400;
        16'hD108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD10C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD110 : rd_rsp_data <= 32'h0100021A;
        16'hD114 : rd_rsp_data <= 32'h00000400;
        16'hD11C : rd_rsp_data <= 32'h00001800;
        16'hD128 : rd_rsp_data <= 32'h00640000;
        16'hD130 : rd_rsp_data <= 32'h00411421;
        16'hD138 : rd_rsp_data <= 32'h00010101;
        16'hD140 : rd_rsp_data <= 32'h0000AA55;
        16'hD144 : rd_rsp_data <= 32'h0000AA55;
        16'hD148 : rd_rsp_data <= 32'h0000AA55;
        16'hD150 : rd_rsp_data <= 32'h01010100;
        16'hD158 : rd_rsp_data <= 32'h80000000;
        16'hD15C : rd_rsp_data <= 32'h80000000;
        16'hD160 : rd_rsp_data <= 32'h80000000;
        16'hD200 : rd_rsp_data <= 32'h01000208;
        16'hD204 : rd_rsp_data <= 32'h00000400;
        16'hD208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD20C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD210 : rd_rsp_data <= 32'h0100021A;
        16'hD214 : rd_rsp_data <= 32'h00000400;
        16'hD21C : rd_rsp_data <= 32'h00001800;
        16'hD228 : rd_rsp_data <= 32'h01040000;
        16'hD230 : rd_rsp_data <= 32'h00411421;
        16'hD238 : rd_rsp_data <= 32'h00010101;
        16'hD240 : rd_rsp_data <= 32'h0000AA55;
        16'hD244 : rd_rsp_data <= 32'h0000AA55;
        16'hD248 : rd_rsp_data <= 32'h0000AA55;
        16'hD250 : rd_rsp_data <= 32'h01010100;
        16'hD258 : rd_rsp_data <= 32'h80000000;
        16'hD25C : rd_rsp_data <= 32'h80000000;
        16'hD260 : rd_rsp_data <= 32'h80000000;
        16'hD300 : rd_rsp_data <= 32'h01000208;
        16'hD304 : rd_rsp_data <= 32'h00000400;
        16'hD308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD30C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD310 : rd_rsp_data <= 32'h0100021A;
        16'hD314 : rd_rsp_data <= 32'h00000400;
        16'hD31C : rd_rsp_data <= 32'h00001800;
        16'hD328 : rd_rsp_data <= 32'h00640000;
        16'hD330 : rd_rsp_data <= 32'h00411421;
        16'hD338 : rd_rsp_data <= 32'h00010101;
        16'hD340 : rd_rsp_data <= 32'h0000AA55;
        16'hD344 : rd_rsp_data <= 32'h0000AA55;
        16'hD348 : rd_rsp_data <= 32'h0000AA55;
        16'hD350 : rd_rsp_data <= 32'h01010100;
        16'hD358 : rd_rsp_data <= 32'h80000000;
        16'hD35C : rd_rsp_data <= 32'h80000000;
        16'hD360 : rd_rsp_data <= 32'h80000000;
        16'hD400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD40C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD41C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD42C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD43C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD44C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD45C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD46C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD47C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD48C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD49C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD4FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD50C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD51C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD52C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD53C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD54C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD55C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD56C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD57C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD58C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD59C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD5FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD60C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD61C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD62C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD63C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD64C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD65C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD66C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD67C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD68C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD69C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD6FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD70C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD71C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD72C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD73C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD74C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD75C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD76C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD77C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD78C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD79C : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD7FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD800 : rd_rsp_data <= 32'h08008001;
        16'hD804 : rd_rsp_data <= 32'h00000100;
        16'hD808 : rd_rsp_data <= 32'h00000100;
        16'hD80C : rd_rsp_data <= 32'hD0000088;
        16'hD810 : rd_rsp_data <= 32'hD0000088;
        16'hD814 : rd_rsp_data <= 32'h00000002;
        16'hD81C : rd_rsp_data <= 32'h00018200;
        16'hD824 : rd_rsp_data <= 32'h130C3200;
        16'hD830 : rd_rsp_data <= 32'h004000AA;
        16'hD834 : rd_rsp_data <= 32'h000004BF;
        16'hD83C : rd_rsp_data <= 32'h00010820;
        16'hD840 : rd_rsp_data <= 32'h8362E297;
        16'hD844 : rd_rsp_data <= 32'h00000012;
        16'hD858 : rd_rsp_data <= 32'h38857E00;
        16'hD85C : rd_rsp_data <= 32'h0000000F;
        16'hD860 : rd_rsp_data <= 32'h00010200;
        16'hD874 : rd_rsp_data <= 32'h00000010;
        16'hD878 : rd_rsp_data <= 32'h00001844;
        16'hD87C : rd_rsp_data <= 32'h00001844;
        16'hD880 : rd_rsp_data <= 32'h24504030;
        16'hD890 : rd_rsp_data <= 32'hFFF00000;
        16'hD894 : rd_rsp_data <= 32'h0000007F;
        16'hD8A0 : rd_rsp_data <= 32'h4886AC7B;
        16'hD8A4 : rd_rsp_data <= 32'h00000003;
        16'hD8A8 : rd_rsp_data <= 32'hF58E67E9;
        16'hD8AC : rd_rsp_data <= 32'h00000023;
        16'hD8BC : rd_rsp_data <= 32'h00100000;
        16'hD930 : rd_rsp_data <= 32'h70B40384;
        16'hD934 : rd_rsp_data <= 32'h0400B05A;
        16'hD938 : rd_rsp_data <= 32'h0000000F;
        16'hD93C : rd_rsp_data <= 32'h00301C1C;
        16'hD954 : rd_rsp_data <= 32'h00300100;
        16'hD958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'hD95C : rd_rsp_data <= 32'h00000001;
        16'hD960 : rd_rsp_data <= 32'h038400E1;
        16'hD964 : rd_rsp_data <= 32'h0000005A;
        16'hD968 : rd_rsp_data <= 32'h0001407D;
        16'hD96C : rd_rsp_data <= 32'h00000001;
        16'hD974 : rd_rsp_data <= 32'h000000C6;
        16'hD9B4 : rd_rsp_data <= 32'h0000001F;
        16'hD9B8 : rd_rsp_data <= 32'h00000107;
        16'hE000 : rd_rsp_data <= 32'h27422027;
        16'hE004 : rd_rsp_data <= 32'h01393075;
        16'hE008 : rd_rsp_data <= 32'h49041828;
        16'hE00C : rd_rsp_data <= 32'h0E0E088C;
        16'hE010 : rd_rsp_data <= 32'h16141212;
        16'hE014 : rd_rsp_data <= 32'h18306C48;
        16'hE018 : rd_rsp_data <= 32'h0E0E081A;
        16'hE01C : rd_rsp_data <= 32'h003FF020;
        16'hE020 : rd_rsp_data <= 32'h19191944;
        16'hE024 : rd_rsp_data <= 32'h19191919;
        16'hE028 : rd_rsp_data <= 32'h80000020;
        16'hE02C : rd_rsp_data <= 32'h4E000200;
        16'hE034 : rd_rsp_data <= 32'h060100B8;
        16'hE038 : rd_rsp_data <= 32'h00000C00;
        16'hE040 : rd_rsp_data <= 32'h000200B8;
        16'hE044 : rd_rsp_data <= 32'h00000200;
        16'hE050 : rd_rsp_data <= 32'h060E8912;
        16'hE054 : rd_rsp_data <= 32'h12068076;
        16'hE068 : rd_rsp_data <= 32'h103B2838;
        16'hE06C : rd_rsp_data <= 32'h16404030;
        16'hE070 : rd_rsp_data <= 32'h26280000;
        16'hE074 : rd_rsp_data <= 32'h00000080;
        16'hE078 : rd_rsp_data <= 32'h00300004;
        16'hE088 : rd_rsp_data <= 32'h8FC00029;
        16'hE08C : rd_rsp_data <= 32'h0C008484;
        16'hE090 : rd_rsp_data <= 32'h0C180810;
        16'hE094 : rd_rsp_data <= 32'h08100408;
        16'hE098 : rd_rsp_data <= 32'h040C0206;
        16'hE0A0 : rd_rsp_data <= 32'hD4CA450A;
        16'hE0A8 : rd_rsp_data <= 32'h02540040;
        16'hE0AC : rd_rsp_data <= 32'h0281284B;
        16'hE0B0 : rd_rsp_data <= 32'h0000000F;
        16'hE0B8 : rd_rsp_data <= 32'h08104426;
        16'hE0C0 : rd_rsp_data <= 32'h00200086;
        16'hE0C4 : rd_rsp_data <= 32'h800308E2;
        16'hE0C8 : rd_rsp_data <= 32'h1C483616;
        16'hE0D0 : rd_rsp_data <= 32'h0000000F;
        16'hE0D4 : rd_rsp_data <= 32'h0E64E893;
        16'hE100 : rd_rsp_data <= 32'h80202028;
        16'hE110 : rd_rsp_data <= 32'h00000056;
        16'hE114 : rd_rsp_data <= 32'h00020611;
        16'hE118 : rd_rsp_data <= 32'hFFF080AE;
        16'hE11C : rd_rsp_data <= 32'h0001B20A;
        16'hE120 : rd_rsp_data <= 32'h000000E0;
        16'hE124 : rd_rsp_data <= 32'h00004000;
        16'hE128 : rd_rsp_data <= 32'h20000000;
        16'hE12C : rd_rsp_data <= 32'h00000007;
        16'hE200 : rd_rsp_data <= 32'h30200884;
        16'hE204 : rd_rsp_data <= 32'h4F3F2F40;
        16'hE208 : rd_rsp_data <= 32'h5E56B731;
        16'hE20C : rd_rsp_data <= 32'h00129024;
        16'hE210 : rd_rsp_data <= 32'h00040844;
        16'hE214 : rd_rsp_data <= 32'hC2C3C1E2;
        16'hE218 : rd_rsp_data <= 32'h1B000036;
        16'hE21C : rd_rsp_data <= 32'h3F001B1B;
        16'hE220 : rd_rsp_data <= 32'h33333838;
        16'hE224 : rd_rsp_data <= 32'h0000007F;
        16'hE3E0 : rd_rsp_data <= 32'h013E9828;
        16'hE3E4 : rd_rsp_data <= 32'h0000508D;
        16'hE3F0 : rd_rsp_data <= 32'hA61DE138;
        16'hE3F4 : rd_rsp_data <= 32'hD0ED45A9;
        16'hE400 : rd_rsp_data <= 32'h11002EC3;
        16'hE404 : rd_rsp_data <= 32'h0000000F;
        16'hE40C : rd_rsp_data <= 32'h00000137;
        16'hE410 : rd_rsp_data <= 32'h00200D05;
        16'hE418 : rd_rsp_data <= 32'h02020202;
        16'hE424 : rd_rsp_data <= 32'h00000001;
        16'hE428 : rd_rsp_data <= 32'h01010101;
        16'hE42C : rd_rsp_data <= 32'h00101020;
        16'hE430 : rd_rsp_data <= 32'h23444688;
        16'hE434 : rd_rsp_data <= 32'h00000008;
        16'hE438 : rd_rsp_data <= 32'h275A7640;
        16'hE43C : rd_rsp_data <= 32'h05FC11C5;
        16'hE440 : rd_rsp_data <= 32'h28000600;
        16'hE444 : rd_rsp_data <= 32'h00004000;
        16'hE448 : rd_rsp_data <= 32'h00013880;
        16'hE44C : rd_rsp_data <= 32'h000004B3;
        16'hE450 : rd_rsp_data <= 32'h00000012;
        16'hE454 : rd_rsp_data <= 32'h00000001;
        16'hE458 : rd_rsp_data <= 32'h00001C00;
        16'hE46C : rd_rsp_data <= 32'h00000101;
        16'hE470 : rd_rsp_data <= 32'h00000101;
        16'hE474 : rd_rsp_data <= 32'h00C96FC8;
        16'hE478 : rd_rsp_data <= 32'h00000003;
        16'hE480 : rd_rsp_data <= 32'h23444688;
        16'hE484 : rd_rsp_data <= 32'h00000009;
        16'hE488 : rd_rsp_data <= 32'h0AC4DC14;
        16'hE494 : rd_rsp_data <= 32'h11311022;
        16'hE498 : rd_rsp_data <= 32'h23444688;
        16'hE49C : rd_rsp_data <= 32'h00000008;
        16'hE4B0 : rd_rsp_data <= 32'h0D9B3E84;
        16'hE4B8 : rd_rsp_data <= 32'h23444688;
        16'hE4BC : rd_rsp_data <= 32'h0000001B;
        16'hE4C0 : rd_rsp_data <= 32'h000002C2;
        16'hE4C4 : rd_rsp_data <= 32'h02000140;
        16'hE4C8 : rd_rsp_data <= 32'h0C078000;
        16'hE4D8 : rd_rsp_data <= 32'h00022000;
        16'hE4FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hE5CC : rd_rsp_data <= 32'h3F000000;
        16'hE5D0 : rd_rsp_data <= 32'hE0400000;
        16'hE5D4 : rd_rsp_data <= 32'h26000400;
        16'hE5E0 : rd_rsp_data <= 32'h00002003;
        16'hE5E4 : rd_rsp_data <= 32'h0000000F;
        16'hE5FC : rd_rsp_data <= 32'h08041000;
        16'hE600 : rd_rsp_data <= 32'h80400000;
        16'hE604 : rd_rsp_data <= 32'h8040010E;
        16'hE608 : rd_rsp_data <= 32'h80400201;
        16'hE60C : rd_rsp_data <= 32'h80400302;
        16'hE610 : rd_rsp_data <= 32'h80400405;
        16'hE614 : rd_rsp_data <= 32'h80400503;
        16'hE618 : rd_rsp_data <= 32'h80400604;
        16'hE61C : rd_rsp_data <= 32'h80400707;
        16'hE620 : rd_rsp_data <= 32'h8480080B;
        16'hE624 : rd_rsp_data <= 32'h8480090C;
        16'hE628 : rd_rsp_data <= 32'h80400A06;
        16'hE62C : rd_rsp_data <= 32'h80400B08;
        16'hE630 : rd_rsp_data <= 32'h80000C00;
        16'hE634 : rd_rsp_data <= 32'h80000D02;
        16'hE638 : rd_rsp_data <= 32'h80000E04;
        16'hE63C : rd_rsp_data <= 32'h80000F05;
        16'hE640 : rd_rsp_data <= 32'h80001006;
        16'hE644 : rd_rsp_data <= 32'h80001108;
        16'hE648 : rd_rsp_data <= 32'h8000120D;
        16'hE64C : rd_rsp_data <= 32'h8000130E;
        16'hE650 : rd_rsp_data <= 32'h80001481;
        16'hE654 : rd_rsp_data <= 32'h80001582;
        16'hE658 : rd_rsp_data <= 32'h80001683;
        16'hE65C : rd_rsp_data <= 32'h80001784;
        16'hE660 : rd_rsp_data <= 32'h80001489;
        16'hE664 : rd_rsp_data <= 32'h8000158A;
        16'hE668 : rd_rsp_data <= 32'h8000168B;
        16'hE66C : rd_rsp_data <= 32'h8000178C;
        16'hE670 : rd_rsp_data <= 32'h80001491;
        16'hE674 : rd_rsp_data <= 32'h80001592;
        16'hE678 : rd_rsp_data <= 32'h80001693;
        16'hE67C : rd_rsp_data <= 32'h80001794;
        16'hE680 : rd_rsp_data <= 32'h80001499;
        16'hE684 : rd_rsp_data <= 32'h8000159A;
        16'hE688 : rd_rsp_data <= 32'h8000169B;
        16'hE68C : rd_rsp_data <= 32'h8000179C;
        16'hE690 : rd_rsp_data <= 32'h800014A1;
        16'hE694 : rd_rsp_data <= 32'h800015A2;
        16'hE698 : rd_rsp_data <= 32'h800016A3;
        16'hE69C : rd_rsp_data <= 32'h800017A4;
        16'hE6A0 : rd_rsp_data <= 32'h800014A9;
        16'hE6A4 : rd_rsp_data <= 32'h800015AA;
        16'hE6A8 : rd_rsp_data <= 32'h800016AB;
        16'hE6AC : rd_rsp_data <= 32'h800017AC;
        16'hE6B0 : rd_rsp_data <= 32'h800014B1;
        16'hE6B4 : rd_rsp_data <= 32'h800015B2;
        16'hE6B8 : rd_rsp_data <= 32'h800016B3;
        16'hE6BC : rd_rsp_data <= 32'h800017B4;
        16'hE6C0 : rd_rsp_data <= 32'h800014B9;
        16'hE6C4 : rd_rsp_data <= 32'h800015BA;
        16'hE6C8 : rd_rsp_data <= 32'h800016BB;
        16'hE6CC : rd_rsp_data <= 32'h800017BC;
        16'hE6D0 : rd_rsp_data <= 32'h800014C1;
        16'hE6D4 : rd_rsp_data <= 32'h800015C2;
        16'hE6D8 : rd_rsp_data <= 32'h800016C3;
        16'hE6DC : rd_rsp_data <= 32'h800017C4;
        16'hE6E0 : rd_rsp_data <= 32'h800014C9;
        16'hE6E4 : rd_rsp_data <= 32'h800015CA;
        16'hE6E8 : rd_rsp_data <= 32'h800016CB;
        16'hE6EC : rd_rsp_data <= 32'h800017CC;
        16'hE6F0 : rd_rsp_data <= 32'h800014D1;
        16'hE6F4 : rd_rsp_data <= 32'h800015D2;
        16'hE6F8 : rd_rsp_data <= 32'h800016D3;
        16'hE6FC : rd_rsp_data <= 32'h800017D4;
        16'hE700 : rd_rsp_data <= 32'h800014D9;
        16'hE704 : rd_rsp_data <= 32'h800015DA;
        16'hE708 : rd_rsp_data <= 32'h800016DB;
        16'hE70C : rd_rsp_data <= 32'h800017DC;
        16'hE710 : rd_rsp_data <= 32'h800014E1;
        16'hE714 : rd_rsp_data <= 32'h800015E2;
        16'hE718 : rd_rsp_data <= 32'h800016E3;
        16'hE71C : rd_rsp_data <= 32'h800017E4;
        16'hE720 : rd_rsp_data <= 32'h800014E9;
        16'hE724 : rd_rsp_data <= 32'h800015EA;
        16'hE728 : rd_rsp_data <= 32'h800016EB;
        16'hE72C : rd_rsp_data <= 32'h800017EC;
        16'hE730 : rd_rsp_data <= 32'h800014F1;
        16'hE734 : rd_rsp_data <= 32'h800015F2;
        16'hE738 : rd_rsp_data <= 32'h800016F3;
        16'hE73C : rd_rsp_data <= 32'h800017F4;
        16'hE740 : rd_rsp_data <= 32'h800014F9;
        16'hE744 : rd_rsp_data <= 32'h800015FA;
        16'hE748 : rd_rsp_data <= 32'h800016FB;
        16'hE74C : rd_rsp_data <= 32'h830017FC;
        16'hE750 : rd_rsp_data <= 32'h80001822;
        16'hE754 : rd_rsp_data <= 32'h80001923;
        16'hE758 : rd_rsp_data <= 32'h80001A24;
        16'hE75C : rd_rsp_data <= 32'h80001B25;
        16'hE760 : rd_rsp_data <= 32'h80001C26;
        16'hE764 : rd_rsp_data <= 32'h80001D27;
        16'hE768 : rd_rsp_data <= 32'h80001E28;
        16'hE76C : rd_rsp_data <= 32'h80001F2D;
        16'hE770 : rd_rsp_data <= 32'hC800200A;
        16'hE774 : rd_rsp_data <= 32'hC8002203;
        16'hE778 : rd_rsp_data <= 32'h8040240F;
        16'hE800 : rd_rsp_data <= 32'h27422027;
        16'hE804 : rd_rsp_data <= 32'h01393075;
        16'hE808 : rd_rsp_data <= 32'h49041828;
        16'hE80C : rd_rsp_data <= 32'h0E0E088C;
        16'hE810 : rd_rsp_data <= 32'h16141212;
        16'hE814 : rd_rsp_data <= 32'h18306C48;
        16'hE818 : rd_rsp_data <= 32'h0E0E081A;
        16'hE81C : rd_rsp_data <= 32'h003FF020;
        16'hE820 : rd_rsp_data <= 32'h1919193F;
        16'hE824 : rd_rsp_data <= 32'h19191919;
        16'hE828 : rd_rsp_data <= 32'h80000020;
        16'hE82C : rd_rsp_data <= 32'h4E000200;
        16'hE834 : rd_rsp_data <= 32'h06010178;
        16'hE838 : rd_rsp_data <= 32'h00000C00;
        16'hE840 : rd_rsp_data <= 32'h000201E8;
        16'hE844 : rd_rsp_data <= 32'h00000200;
        16'hE850 : rd_rsp_data <= 32'h060E8912;
        16'hE854 : rd_rsp_data <= 32'h12068076;
        16'hE868 : rd_rsp_data <= 32'h103B2838;
        16'hE86C : rd_rsp_data <= 32'h16404030;
        16'hE870 : rd_rsp_data <= 32'h26280000;
        16'hE874 : rd_rsp_data <= 32'h00000080;
        16'hE878 : rd_rsp_data <= 32'h00300004;
        16'hE888 : rd_rsp_data <= 32'h8FC00029;
        16'hE88C : rd_rsp_data <= 32'h0C008484;
        16'hE890 : rd_rsp_data <= 32'h0C180810;
        16'hE894 : rd_rsp_data <= 32'h08100408;
        16'hE898 : rd_rsp_data <= 32'h040C0206;
        16'hE8A0 : rd_rsp_data <= 32'hD4CA450A;
        16'hE8A8 : rd_rsp_data <= 32'h02540040;
        16'hE8AC : rd_rsp_data <= 32'h0281284B;
        16'hE8B0 : rd_rsp_data <= 32'h0000000F;
        16'hE8B8 : rd_rsp_data <= 32'h08104426;
        16'hE8C0 : rd_rsp_data <= 32'h00200086;
        16'hE8C4 : rd_rsp_data <= 32'h800308E2;
        16'hE8C8 : rd_rsp_data <= 32'h1C483616;
        16'hE8D0 : rd_rsp_data <= 32'h0000000F;
        16'hE8D4 : rd_rsp_data <= 32'h0E64E893;
        16'hE900 : rd_rsp_data <= 32'h80202028;
        16'hE910 : rd_rsp_data <= 32'h00000056;
        16'hE914 : rd_rsp_data <= 32'h00020611;
        16'hE918 : rd_rsp_data <= 32'hFFF080AE;
        16'hE91C : rd_rsp_data <= 32'h0001B20A;
        16'hE920 : rd_rsp_data <= 32'h000000E0;
        16'hE924 : rd_rsp_data <= 32'h00004000;
        16'hE928 : rd_rsp_data <= 32'h20000000;
        16'hE92C : rd_rsp_data <= 32'h00000007;
        16'hEA00 : rd_rsp_data <= 32'h30200884;
        16'hEA04 : rd_rsp_data <= 32'h4F3F2F40;
        16'hEA08 : rd_rsp_data <= 32'h5E56B734;
        16'hEA0C : rd_rsp_data <= 32'h00129024;
        16'hEA10 : rd_rsp_data <= 32'h00040844;
        16'hEA14 : rd_rsp_data <= 32'hC1C5C2DD;
        16'hEA18 : rd_rsp_data <= 32'h1B000036;
        16'hEA1C : rd_rsp_data <= 32'h3F001B1B;
        16'hEA20 : rd_rsp_data <= 32'h33333A3A;
        16'hEA24 : rd_rsp_data <= 32'h0000007F;
        16'hEBE0 : rd_rsp_data <= 32'h013E9828;
        16'hEBE4 : rd_rsp_data <= 32'h0000508D;
        16'hEBF0 : rd_rsp_data <= 32'h1DCA318B;
        16'hEBF4 : rd_rsp_data <= 32'h864C9844;
        16'hEC00 : rd_rsp_data <= 32'h11002EC3;
        16'hEC04 : rd_rsp_data <= 32'h0000000F;
        16'hEC0C : rd_rsp_data <= 32'h00000137;
        16'hEC10 : rd_rsp_data <= 32'h00200D05;
        16'hEC18 : rd_rsp_data <= 32'h02020202;
        16'hEC24 : rd_rsp_data <= 32'h00000001;
        16'hEC28 : rd_rsp_data <= 32'h01010101;
        16'hEC2C : rd_rsp_data <= 32'h00101020;
        16'hEC30 : rd_rsp_data <= 32'h23444688;
        16'hEC34 : rd_rsp_data <= 32'h00000008;
        16'hEC38 : rd_rsp_data <= 32'h275A7640;
        16'hEC3C : rd_rsp_data <= 32'h05FC11C5;
        16'hEC40 : rd_rsp_data <= 32'h28000600;
        16'hEC44 : rd_rsp_data <= 32'h00004000;
        16'hEC48 : rd_rsp_data <= 32'h00013880;
        16'hEC4C : rd_rsp_data <= 32'h000004B3;
        16'hEC50 : rd_rsp_data <= 32'h00000012;
        16'hEC54 : rd_rsp_data <= 32'h00000001;
        16'hEC58 : rd_rsp_data <= 32'h00001C00;
        16'hEC6C : rd_rsp_data <= 32'h00000101;
        16'hEC70 : rd_rsp_data <= 32'h00000101;
        16'hEC74 : rd_rsp_data <= 32'h00FF3948;
        16'hEC78 : rd_rsp_data <= 32'h00000004;
        16'hEC80 : rd_rsp_data <= 32'h23444688;
        16'hEC88 : rd_rsp_data <= 32'h0AC4DC14;
        16'hEC94 : rd_rsp_data <= 32'h11311022;
        16'hEC98 : rd_rsp_data <= 32'h23444688;
        16'hEC9C : rd_rsp_data <= 32'h00000008;
        16'hECB0 : rd_rsp_data <= 32'h0D9B43BB;
        16'hECB8 : rd_rsp_data <= 32'h23444688;
        16'hECBC : rd_rsp_data <= 32'h00000012;
        16'hECC0 : rd_rsp_data <= 32'h000002C2;
        16'hECC4 : rd_rsp_data <= 32'h02000140;
        16'hECC8 : rd_rsp_data <= 32'h0C078000;
        16'hECD8 : rd_rsp_data <= 32'h09BA6FD6;
        16'hECDC : rd_rsp_data <= 32'hD43F083F;
        16'hECFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hEDCC : rd_rsp_data <= 32'h3F000000;
        16'hEDD0 : rd_rsp_data <= 32'hE0400000;
        16'hEDD4 : rd_rsp_data <= 32'h26000400;
        16'hEDE0 : rd_rsp_data <= 32'h00002003;
        16'hEDE4 : rd_rsp_data <= 32'h0000000F;
        16'hEDFC : rd_rsp_data <= 32'h08041000;
        16'hEE00 : rd_rsp_data <= 32'h80400000;
        16'hEE04 : rd_rsp_data <= 32'h8040010E;
        16'hEE08 : rd_rsp_data <= 32'h80400201;
        16'hEE0C : rd_rsp_data <= 32'h80400302;
        16'hEE10 : rd_rsp_data <= 32'h80400405;
        16'hEE14 : rd_rsp_data <= 32'h80400503;
        16'hEE18 : rd_rsp_data <= 32'h80400604;
        16'hEE1C : rd_rsp_data <= 32'h80400707;
        16'hEE20 : rd_rsp_data <= 32'h8480080B;
        16'hEE24 : rd_rsp_data <= 32'h8480090C;
        16'hEE28 : rd_rsp_data <= 32'h80400A06;
        16'hEE2C : rd_rsp_data <= 32'h80400B08;
        16'hEE30 : rd_rsp_data <= 32'h80000C00;
        16'hEE34 : rd_rsp_data <= 32'h80000D02;
        16'hEE38 : rd_rsp_data <= 32'h80000E04;
        16'hEE3C : rd_rsp_data <= 32'h80000F05;
        16'hEE40 : rd_rsp_data <= 32'h80001006;
        16'hEE44 : rd_rsp_data <= 32'h80001108;
        16'hEE48 : rd_rsp_data <= 32'h8000120D;
        16'hEE4C : rd_rsp_data <= 32'h8000130E;
        16'hEE50 : rd_rsp_data <= 32'h80001481;
        16'hEE54 : rd_rsp_data <= 32'h80001582;
        16'hEE58 : rd_rsp_data <= 32'h80001683;
        16'hEE5C : rd_rsp_data <= 32'h80001784;
        16'hEE60 : rd_rsp_data <= 32'h80001489;
        16'hEE64 : rd_rsp_data <= 32'h8000158A;
        16'hEE68 : rd_rsp_data <= 32'h8000168B;
        16'hEE6C : rd_rsp_data <= 32'h8000178C;
        16'hEE70 : rd_rsp_data <= 32'h80001491;
        16'hEE74 : rd_rsp_data <= 32'h80001592;
        16'hEE78 : rd_rsp_data <= 32'h80001693;
        16'hEE7C : rd_rsp_data <= 32'h80001794;
        16'hEE80 : rd_rsp_data <= 32'h80001499;
        16'hEE84 : rd_rsp_data <= 32'h8000159A;
        16'hEE88 : rd_rsp_data <= 32'h8000169B;
        16'hEE8C : rd_rsp_data <= 32'h8000179C;
        16'hEE90 : rd_rsp_data <= 32'h800014A1;
        16'hEE94 : rd_rsp_data <= 32'h800015A2;
        16'hEE98 : rd_rsp_data <= 32'h800016A3;
        16'hEE9C : rd_rsp_data <= 32'h800017A4;
        16'hEEA0 : rd_rsp_data <= 32'h800014A9;
        16'hEEA4 : rd_rsp_data <= 32'h800015AA;
        16'hEEA8 : rd_rsp_data <= 32'h800016AB;
        16'hEEAC : rd_rsp_data <= 32'h800017AC;
        16'hEEB0 : rd_rsp_data <= 32'h800014B1;
        16'hEEB4 : rd_rsp_data <= 32'h800015B2;
        16'hEEB8 : rd_rsp_data <= 32'h800016B3;
        16'hEEBC : rd_rsp_data <= 32'h800017B4;
        16'hEEC0 : rd_rsp_data <= 32'h800014B9;
        16'hEEC4 : rd_rsp_data <= 32'h800015BA;
        16'hEEC8 : rd_rsp_data <= 32'h800016BB;
        16'hEECC : rd_rsp_data <= 32'h800017BC;
        16'hEED0 : rd_rsp_data <= 32'h800014C1;
        16'hEED4 : rd_rsp_data <= 32'h800015C2;
        16'hEED8 : rd_rsp_data <= 32'h800016C3;
        16'hEEDC : rd_rsp_data <= 32'h800017C4;
        16'hEEE0 : rd_rsp_data <= 32'h800014C9;
        16'hEEE4 : rd_rsp_data <= 32'h800015CA;
        16'hEEE8 : rd_rsp_data <= 32'h800016CB;
        16'hEEEC : rd_rsp_data <= 32'h800017CC;
        16'hEEF0 : rd_rsp_data <= 32'h800014D1;
        16'hEEF4 : rd_rsp_data <= 32'h800015D2;
        16'hEEF8 : rd_rsp_data <= 32'h800016D3;
        16'hEEFC : rd_rsp_data <= 32'h800017D4;
        16'hEF00 : rd_rsp_data <= 32'h800014D9;
        16'hEF04 : rd_rsp_data <= 32'h800015DA;
        16'hEF08 : rd_rsp_data <= 32'h800016DB;
        16'hEF0C : rd_rsp_data <= 32'h800017DC;
        16'hEF10 : rd_rsp_data <= 32'h800014E1;
        16'hEF14 : rd_rsp_data <= 32'h800015E2;
        16'hEF18 : rd_rsp_data <= 32'h800016E3;
        16'hEF1C : rd_rsp_data <= 32'h800017E4;
        16'hEF20 : rd_rsp_data <= 32'h800014E9;
        16'hEF24 : rd_rsp_data <= 32'h800015EA;
        16'hEF28 : rd_rsp_data <= 32'h800016EB;
        16'hEF2C : rd_rsp_data <= 32'h800017EC;
        16'hEF30 : rd_rsp_data <= 32'h800014F1;
        16'hEF34 : rd_rsp_data <= 32'h800015F2;
        16'hEF38 : rd_rsp_data <= 32'h800016F3;
        16'hEF3C : rd_rsp_data <= 32'h800017F4;
        16'hEF40 : rd_rsp_data <= 32'h800014F9;
        16'hEF44 : rd_rsp_data <= 32'h800015FA;
        16'hEF48 : rd_rsp_data <= 32'h800016FB;
        16'hEF4C : rd_rsp_data <= 32'h830017FC;
        16'hEF50 : rd_rsp_data <= 32'h80001822;
        16'hEF54 : rd_rsp_data <= 32'h80001923;
        16'hEF58 : rd_rsp_data <= 32'h80001A24;
        16'hEF5C : rd_rsp_data <= 32'h80001B25;
        16'hEF60 : rd_rsp_data <= 32'h80001C26;
        16'hEF64 : rd_rsp_data <= 32'h80001D27;
        16'hEF68 : rd_rsp_data <= 32'h80001E28;
        16'hEF6C : rd_rsp_data <= 32'h80001F2D;
        16'hEF70 : rd_rsp_data <= 32'hC800200A;
        16'hEF74 : rd_rsp_data <= 32'hC8002203;
        16'hEF78 : rd_rsp_data <= 32'h8040240F;
        16'hF000 : rd_rsp_data <= 32'h27422027;
        16'hF004 : rd_rsp_data <= 32'h01393075;
        16'hF008 : rd_rsp_data <= 32'h49041828;
        16'hF00C : rd_rsp_data <= 32'h0E0E088C;
        16'hF010 : rd_rsp_data <= 32'h16141212;
        16'hF014 : rd_rsp_data <= 32'h18306C48;
        16'hF018 : rd_rsp_data <= 32'h0E0E081A;
        16'hF01C : rd_rsp_data <= 32'h003FF020;
        16'hF020 : rd_rsp_data <= 32'h19191944;
        16'hF024 : rd_rsp_data <= 32'h19191919;
        16'hF028 : rd_rsp_data <= 32'h80000020;
        16'hF02C : rd_rsp_data <= 32'h4E000200;
        16'hF034 : rd_rsp_data <= 32'h06010118;
        16'hF038 : rd_rsp_data <= 32'h00000C00;
        16'hF040 : rd_rsp_data <= 32'h00020118;
        16'hF044 : rd_rsp_data <= 32'h00000200;
        16'hF050 : rd_rsp_data <= 32'h060E8912;
        16'hF054 : rd_rsp_data <= 32'h12068076;
        16'hF068 : rd_rsp_data <= 32'h103B2838;
        16'hF06C : rd_rsp_data <= 32'h16404030;
        16'hF070 : rd_rsp_data <= 32'h26280000;
        16'hF074 : rd_rsp_data <= 32'h00000080;
        16'hF078 : rd_rsp_data <= 32'h00300004;
        16'hF088 : rd_rsp_data <= 32'h8FC00029;
        16'hF08C : rd_rsp_data <= 32'h0C008484;
        16'hF090 : rd_rsp_data <= 32'h0C180810;
        16'hF094 : rd_rsp_data <= 32'h08100408;
        16'hF098 : rd_rsp_data <= 32'h040C0206;
        16'hF0A0 : rd_rsp_data <= 32'hD4CA450A;
        16'hF0A8 : rd_rsp_data <= 32'h02540040;
        16'hF0AC : rd_rsp_data <= 32'h0281284B;
        16'hF0B0 : rd_rsp_data <= 32'h0000000F;
        16'hF0B8 : rd_rsp_data <= 32'h08104426;
        16'hF0C0 : rd_rsp_data <= 32'h00200086;
        16'hF0C4 : rd_rsp_data <= 32'h800308E2;
        16'hF0C8 : rd_rsp_data <= 32'h1C483616;
        16'hF0D0 : rd_rsp_data <= 32'h0000000F;
        16'hF0D4 : rd_rsp_data <= 32'h0E64E893;
        16'hF100 : rd_rsp_data <= 32'h80202028;
        16'hF110 : rd_rsp_data <= 32'h00000056;
        16'hF114 : rd_rsp_data <= 32'h00020611;
        16'hF118 : rd_rsp_data <= 32'hFFF080AE;
        16'hF11C : rd_rsp_data <= 32'h0001B20A;
        16'hF120 : rd_rsp_data <= 32'h000000E0;
        16'hF124 : rd_rsp_data <= 32'h00004000;
        16'hF128 : rd_rsp_data <= 32'h20000000;
        16'hF12C : rd_rsp_data <= 32'h00000007;
        16'hF200 : rd_rsp_data <= 32'h30200884;
        16'hF204 : rd_rsp_data <= 32'h4F3F2F40;
        16'hF208 : rd_rsp_data <= 32'h5E56B731;
        16'hF20C : rd_rsp_data <= 32'h00129024;
        16'hF210 : rd_rsp_data <= 32'h00040844;
        16'hF214 : rd_rsp_data <= 32'hC2C3C1E2;
        16'hF218 : rd_rsp_data <= 32'h1B000036;
        16'hF21C : rd_rsp_data <= 32'h3F001B1B;
        16'hF220 : rd_rsp_data <= 32'h33333838;
        16'hF224 : rd_rsp_data <= 32'h0000007F;
        16'hF3E0 : rd_rsp_data <= 32'h013E9828;
        16'hF3E4 : rd_rsp_data <= 32'h0000508D;
        16'hF3F0 : rd_rsp_data <= 32'h919B9E0F;
        16'hF3F4 : rd_rsp_data <= 32'hEBAD8D1B;
        16'hF400 : rd_rsp_data <= 32'h11002EC3;
        16'hF404 : rd_rsp_data <= 32'h0000000F;
        16'hF40C : rd_rsp_data <= 32'h00000137;
        16'hF410 : rd_rsp_data <= 32'h00200D05;
        16'hF418 : rd_rsp_data <= 32'h02020202;
        16'hF424 : rd_rsp_data <= 32'h00000001;
        16'hF428 : rd_rsp_data <= 32'h01010101;
        16'hF42C : rd_rsp_data <= 32'h00101020;
        16'hF430 : rd_rsp_data <= 32'h23444688;
        16'hF434 : rd_rsp_data <= 32'h00000008;
        16'hF438 : rd_rsp_data <= 32'h275A7640;
        16'hF43C : rd_rsp_data <= 32'h05FC11C5;
        16'hF440 : rd_rsp_data <= 32'h28000600;
        16'hF444 : rd_rsp_data <= 32'h00004000;
        16'hF448 : rd_rsp_data <= 32'h00013880;
        16'hF44C : rd_rsp_data <= 32'h000004B3;
        16'hF450 : rd_rsp_data <= 32'h00000012;
        16'hF454 : rd_rsp_data <= 32'h00000001;
        16'hF458 : rd_rsp_data <= 32'h00001C00;
        16'hF46C : rd_rsp_data <= 32'h00000101;
        16'hF470 : rd_rsp_data <= 32'h00000101;
        16'hF474 : rd_rsp_data <= 32'h00C96FC8;
        16'hF478 : rd_rsp_data <= 32'h00000003;
        16'hF480 : rd_rsp_data <= 32'h23444688;
        16'hF484 : rd_rsp_data <= 32'h00000009;
        16'hF488 : rd_rsp_data <= 32'h0AC4DC14;
        16'hF494 : rd_rsp_data <= 32'h11311022;
        16'hF498 : rd_rsp_data <= 32'h23444688;
        16'hF49C : rd_rsp_data <= 32'h00000008;
        16'hF4B0 : rd_rsp_data <= 32'h0D9B3E84;
        16'hF4B8 : rd_rsp_data <= 32'h23444688;
        16'hF4BC : rd_rsp_data <= 32'h0000001B;
        16'hF4C0 : rd_rsp_data <= 32'h000002C2;
        16'hF4C4 : rd_rsp_data <= 32'h02000140;
        16'hF4C8 : rd_rsp_data <= 32'h0C078000;
        16'hF4D8 : rd_rsp_data <= 32'h00022000;
        16'hF4FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'hF5CC : rd_rsp_data <= 32'h3F000000;
        16'hF5D0 : rd_rsp_data <= 32'hE0400000;
        16'hF5D4 : rd_rsp_data <= 32'h26000400;
        16'hF5E0 : rd_rsp_data <= 32'h00002003;
        16'hF5E4 : rd_rsp_data <= 32'h0000000F;
        16'hF5FC : rd_rsp_data <= 32'h08041000;
        16'hF600 : rd_rsp_data <= 32'h80400000;
        16'hF604 : rd_rsp_data <= 32'h8040010E;
        16'hF608 : rd_rsp_data <= 32'h80400201;
        16'hF60C : rd_rsp_data <= 32'h80400302;
        16'hF610 : rd_rsp_data <= 32'h80400405;
        16'hF614 : rd_rsp_data <= 32'h80400503;
        16'hF618 : rd_rsp_data <= 32'h80400604;
        16'hF61C : rd_rsp_data <= 32'h80400707;
        16'hF620 : rd_rsp_data <= 32'h8480080B;
        16'hF624 : rd_rsp_data <= 32'h8480090C;
        16'hF628 : rd_rsp_data <= 32'h80400A06;
        16'hF62C : rd_rsp_data <= 32'h80400B08;
        16'hF630 : rd_rsp_data <= 32'h80000C00;
        16'hF634 : rd_rsp_data <= 32'h80000D02;
        16'hF638 : rd_rsp_data <= 32'h80000E04;
        16'hF63C : rd_rsp_data <= 32'h80000F05;
        16'hF640 : rd_rsp_data <= 32'h80001006;
        16'hF644 : rd_rsp_data <= 32'h80001108;
        16'hF648 : rd_rsp_data <= 32'h8000120D;
        16'hF64C : rd_rsp_data <= 32'h8000130E;
        16'hF650 : rd_rsp_data <= 32'h80001481;
        16'hF654 : rd_rsp_data <= 32'h80001582;
        16'hF658 : rd_rsp_data <= 32'h80001683;
        16'hF65C : rd_rsp_data <= 32'h80001784;
        16'hF660 : rd_rsp_data <= 32'h80001489;
        16'hF664 : rd_rsp_data <= 32'h8000158A;
        16'hF668 : rd_rsp_data <= 32'h8000168B;
        16'hF66C : rd_rsp_data <= 32'h8000178C;
        16'hF670 : rd_rsp_data <= 32'h80001491;
        16'hF674 : rd_rsp_data <= 32'h80001592;
        16'hF678 : rd_rsp_data <= 32'h80001693;
        16'hF67C : rd_rsp_data <= 32'h80001794;
        16'hF680 : rd_rsp_data <= 32'h80001499;
        16'hF684 : rd_rsp_data <= 32'h8000159A;
        16'hF688 : rd_rsp_data <= 32'h8000169B;
        16'hF68C : rd_rsp_data <= 32'h8000179C;
        16'hF690 : rd_rsp_data <= 32'h800014A1;
        16'hF694 : rd_rsp_data <= 32'h800015A2;
        16'hF698 : rd_rsp_data <= 32'h800016A3;
        16'hF69C : rd_rsp_data <= 32'h800017A4;
        16'hF6A0 : rd_rsp_data <= 32'h800014A9;
        16'hF6A4 : rd_rsp_data <= 32'h800015AA;
        16'hF6A8 : rd_rsp_data <= 32'h800016AB;
        16'hF6AC : rd_rsp_data <= 32'h800017AC;
        16'hF6B0 : rd_rsp_data <= 32'h800014B1;
        16'hF6B4 : rd_rsp_data <= 32'h800015B2;
        16'hF6B8 : rd_rsp_data <= 32'h800016B3;
        16'hF6BC : rd_rsp_data <= 32'h800017B4;
        16'hF6C0 : rd_rsp_data <= 32'h800014B9;
        16'hF6C4 : rd_rsp_data <= 32'h800015BA;
        16'hF6C8 : rd_rsp_data <= 32'h800016BB;
        16'hF6CC : rd_rsp_data <= 32'h800017BC;
        16'hF6D0 : rd_rsp_data <= 32'h800014C1;
        16'hF6D4 : rd_rsp_data <= 32'h800015C2;
        16'hF6D8 : rd_rsp_data <= 32'h800016C3;
        16'hF6DC : rd_rsp_data <= 32'h800017C4;
        16'hF6E0 : rd_rsp_data <= 32'h800014C9;
        16'hF6E4 : rd_rsp_data <= 32'h800015CA;
        16'hF6E8 : rd_rsp_data <= 32'h800016CB;
        16'hF6EC : rd_rsp_data <= 32'h800017CC;
        16'hF6F0 : rd_rsp_data <= 32'h800014D1;
        16'hF6F4 : rd_rsp_data <= 32'h800015D2;
        16'hF6F8 : rd_rsp_data <= 32'h800016D3;
        16'hF6FC : rd_rsp_data <= 32'h800017D4;
        16'hF700 : rd_rsp_data <= 32'h800014D9;
        16'hF704 : rd_rsp_data <= 32'h800015DA;
        16'hF708 : rd_rsp_data <= 32'h800016DB;
        16'hF70C : rd_rsp_data <= 32'h800017DC;
        16'hF710 : rd_rsp_data <= 32'h800014E1;
        16'hF714 : rd_rsp_data <= 32'h800015E2;
        16'hF718 : rd_rsp_data <= 32'h800016E3;
        16'hF71C : rd_rsp_data <= 32'h800017E4;
        16'hF720 : rd_rsp_data <= 32'h800014E9;
        16'hF724 : rd_rsp_data <= 32'h800015EA;
        16'hF728 : rd_rsp_data <= 32'h800016EB;
        16'hF72C : rd_rsp_data <= 32'h800017EC;
        16'hF730 : rd_rsp_data <= 32'h800014F1;
        16'hF734 : rd_rsp_data <= 32'h800015F2;
        16'hF738 : rd_rsp_data <= 32'h800016F3;
        16'hF73C : rd_rsp_data <= 32'h800017F4;
        16'hF740 : rd_rsp_data <= 32'h800014F9;
        16'hF744 : rd_rsp_data <= 32'h800015FA;
        16'hF748 : rd_rsp_data <= 32'h800016FB;
        16'hF74C : rd_rsp_data <= 32'h830017FC;
        16'hF750 : rd_rsp_data <= 32'h80001822;
        16'hF754 : rd_rsp_data <= 32'h80001923;
        16'hF758 : rd_rsp_data <= 32'h80001A24;
        16'hF75C : rd_rsp_data <= 32'h80001B25;
        16'hF760 : rd_rsp_data <= 32'h80001C26;
        16'hF764 : rd_rsp_data <= 32'h80001D27;
        16'hF768 : rd_rsp_data <= 32'h80001E28;
        16'hF76C : rd_rsp_data <= 32'h80001F2D;
        16'hF770 : rd_rsp_data <= 32'hC800200A;
        16'hF774 : rd_rsp_data <= 32'hC8002203;
        16'hF778 : rd_rsp_data <= 32'h8040240F;
        16'h10000 : rd_rsp_data <= 32'h01010208;
        16'h10004 : rd_rsp_data <= 32'h00000400;
        16'h10008 : rd_rsp_data <= 32'h4101861F;
        16'h1000C : rd_rsp_data <= 32'h00001408;
        16'h10010 : rd_rsp_data <= 32'h01000208;
        16'h10014 : rd_rsp_data <= 32'h00000400;
        16'h10018 : rd_rsp_data <= 32'h0100021A;
        16'h1001C : rd_rsp_data <= 32'h00000400;
        16'h10020 : rd_rsp_data <= 32'h01000208;
        16'h10024 : rd_rsp_data <= 32'h00000400;
        16'h10028 : rd_rsp_data <= 32'h01000608;
        16'h1002C : rd_rsp_data <= 32'h00001500;
        16'h10030 : rd_rsp_data <= 32'h01000208;
        16'h10034 : rd_rsp_data <= 32'h00000400;
        16'h10038 : rd_rsp_data <= 32'h0100020A;
        16'h1003C : rd_rsp_data <= 32'h00000400;
        16'h10040 : rd_rsp_data <= 32'h0100020A;
        16'h10044 : rd_rsp_data <= 32'h00000400;
        16'h10068 : rd_rsp_data <= 32'h00000010;
        16'h10100 : rd_rsp_data <= 32'h000000FE;
        16'h10120 : rd_rsp_data <= 32'h00FFFFFF;
        16'h1012C : rd_rsp_data <= 32'h00000B63;
        16'h10130 : rd_rsp_data <= 32'h0000000C;
        16'h10150 : rd_rsp_data <= 32'h00000001;
        16'h10170 : rd_rsp_data <= 32'h00001FF7;
        16'h1017C : rd_rsp_data <= 32'h00000004;
        16'h10180 : rd_rsp_data <= 32'hAD7FFFFF;
        16'h10184 : rd_rsp_data <= 32'h00000004;
        16'h10188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10190 : rd_rsp_data <= 32'h00010000;
        16'h10198 : rd_rsp_data <= 32'h03082404;
        16'h10200 : rd_rsp_data <= 32'h0011C000;
        16'h10204 : rd_rsp_data <= 32'hFFFFC000;
        16'h10208 : rd_rsp_data <= 32'h01010210;
        16'h1020C : rd_rsp_data <= 32'h00000400;
        16'h10210 : rd_rsp_data <= 32'h01010210;
        16'h10214 : rd_rsp_data <= 32'h00000400;
        16'h10218 : rd_rsp_data <= 32'h01010210;
        16'h1021C : rd_rsp_data <= 32'h00000400;
        16'h10228 : rd_rsp_data <= 32'h01010210;
        16'h1022C : rd_rsp_data <= 32'h00000400;
        16'h10230 : rd_rsp_data <= 32'h01010210;
        16'h10234 : rd_rsp_data <= 32'h00000400;
        16'h10238 : rd_rsp_data <= 32'h01010210;
        16'h1023C : rd_rsp_data <= 32'h00000400;
        16'h10240 : rd_rsp_data <= 32'h00120000;
        16'h10244 : rd_rsp_data <= 32'hFFFFC000;
        16'h10248 : rd_rsp_data <= 32'h01010210;
        16'h1024C : rd_rsp_data <= 32'h00000400;
        16'h10250 : rd_rsp_data <= 32'h01010210;
        16'h10254 : rd_rsp_data <= 32'h00020400;
        16'h10258 : rd_rsp_data <= 32'h01010210;
        16'h1025C : rd_rsp_data <= 32'h00020400;
        16'h10268 : rd_rsp_data <= 32'h01010210;
        16'h1026C : rd_rsp_data <= 32'h00000400;
        16'h10270 : rd_rsp_data <= 32'h01010210;
        16'h10274 : rd_rsp_data <= 32'h00000400;
        16'h10278 : rd_rsp_data <= 32'h01010210;
        16'h1027C : rd_rsp_data <= 32'h00000400;
        16'h10288 : rd_rsp_data <= 32'h01010210;
        16'h1028C : rd_rsp_data <= 32'h00000400;
        16'h10290 : rd_rsp_data <= 32'h01010210;
        16'h10294 : rd_rsp_data <= 32'h00000400;
        16'h10298 : rd_rsp_data <= 32'h01010210;
        16'h1029C : rd_rsp_data <= 32'h00000400;
        16'h102A8 : rd_rsp_data <= 32'h01010210;
        16'h102AC : rd_rsp_data <= 32'h00000400;
        16'h102B0 : rd_rsp_data <= 32'h01010210;
        16'h102B4 : rd_rsp_data <= 32'h00000400;
        16'h102B8 : rd_rsp_data <= 32'h01010210;
        16'h102BC : rd_rsp_data <= 32'h00000400;
        16'h102C8 : rd_rsp_data <= 32'h01010210;
        16'h102CC : rd_rsp_data <= 32'h00000400;
        16'h102D0 : rd_rsp_data <= 32'h01010210;
        16'h102D4 : rd_rsp_data <= 32'h00000400;
        16'h102D8 : rd_rsp_data <= 32'h01010210;
        16'h102DC : rd_rsp_data <= 32'h00000400;
        16'h102E8 : rd_rsp_data <= 32'h01010210;
        16'h102EC : rd_rsp_data <= 32'h00000400;
        16'h102F0 : rd_rsp_data <= 32'h01010210;
        16'h102F4 : rd_rsp_data <= 32'h00000400;
        16'h102F8 : rd_rsp_data <= 32'h01010210;
        16'h102FC : rd_rsp_data <= 32'h00000400;
        16'h10300 : rd_rsp_data <= 32'h00124000;
        16'h10304 : rd_rsp_data <= 32'hFFFFF000;
        16'h10308 : rd_rsp_data <= 32'h01010210;
        16'h1030C : rd_rsp_data <= 32'h00000400;
        16'h10310 : rd_rsp_data <= 32'h01000210;
        16'h10314 : rd_rsp_data <= 32'h02000400;
        16'h10318 : rd_rsp_data <= 32'h01000210;
        16'h1031C : rd_rsp_data <= 32'h02000400;
        16'h10328 : rd_rsp_data <= 32'h01010210;
        16'h1032C : rd_rsp_data <= 32'h00000400;
        16'h10330 : rd_rsp_data <= 32'h01010210;
        16'h10334 : rd_rsp_data <= 32'h00000400;
        16'h10338 : rd_rsp_data <= 32'h01010210;
        16'h1033C : rd_rsp_data <= 32'h00000400;
        16'h10348 : rd_rsp_data <= 32'h01010210;
        16'h1034C : rd_rsp_data <= 32'h00000400;
        16'h10350 : rd_rsp_data <= 32'h01010210;
        16'h10354 : rd_rsp_data <= 32'h00000400;
        16'h10358 : rd_rsp_data <= 32'h01010210;
        16'h1035C : rd_rsp_data <= 32'h00000400;
        16'h10368 : rd_rsp_data <= 32'h01010210;
        16'h1036C : rd_rsp_data <= 32'h00000400;
        16'h10370 : rd_rsp_data <= 32'h01010210;
        16'h10374 : rd_rsp_data <= 32'h00000400;
        16'h10378 : rd_rsp_data <= 32'h01010210;
        16'h1037C : rd_rsp_data <= 32'h00000400;
        16'h10380 : rd_rsp_data <= 32'h00125000;
        16'h10384 : rd_rsp_data <= 32'hFFFFFFE0;
        16'h10388 : rd_rsp_data <= 32'h01010210;
        16'h1038C : rd_rsp_data <= 32'h00000400;
        16'h10390 : rd_rsp_data <= 32'h01010210;
        16'h10394 : rd_rsp_data <= 32'h00000400;
        16'h10398 : rd_rsp_data <= 32'h01010210;
        16'h1039C : rd_rsp_data <= 32'h00000400;
        16'h103A8 : rd_rsp_data <= 32'h01000200;
        16'h103AC : rd_rsp_data <= 32'h00000400;
        16'h103C0 : rd_rsp_data <= 32'h00125020;
        16'h103C4 : rd_rsp_data <= 32'hFFFFFFE0;
        16'h103C8 : rd_rsp_data <= 32'h01010210;
        16'h103CC : rd_rsp_data <= 32'h00000400;
        16'h103D0 : rd_rsp_data <= 32'h01010210;
        16'h103D4 : rd_rsp_data <= 32'h00000400;
        16'h103D8 : rd_rsp_data <= 32'h01010210;
        16'h103DC : rd_rsp_data <= 32'h00000400;
        16'h103E8 : rd_rsp_data <= 32'h01010210;
        16'h103EC : rd_rsp_data <= 32'h00000400;
        16'h103F0 : rd_rsp_data <= 32'h01010210;
        16'h103F4 : rd_rsp_data <= 32'h00000400;
        16'h103F8 : rd_rsp_data <= 32'h01010210;
        16'h103FC : rd_rsp_data <= 32'h00000400;
        16'h10408 : rd_rsp_data <= 32'h01010210;
        16'h1040C : rd_rsp_data <= 32'h00000400;
        16'h10410 : rd_rsp_data <= 32'h01010210;
        16'h10414 : rd_rsp_data <= 32'h00000400;
        16'h10418 : rd_rsp_data <= 32'h01010210;
        16'h1041C : rd_rsp_data <= 32'h00000400;
        16'h10428 : rd_rsp_data <= 32'h01010210;
        16'h1042C : rd_rsp_data <= 32'h00000400;
        16'h10430 : rd_rsp_data <= 32'h01010210;
        16'h10434 : rd_rsp_data <= 32'h00000400;
        16'h10438 : rd_rsp_data <= 32'h01010210;
        16'h1043C : rd_rsp_data <= 32'h00000400;
        16'h10448 : rd_rsp_data <= 32'h01010210;
        16'h1044C : rd_rsp_data <= 32'h00000400;
        16'h10450 : rd_rsp_data <= 32'h01010210;
        16'h10454 : rd_rsp_data <= 32'h00000400;
        16'h10458 : rd_rsp_data <= 32'h01010210;
        16'h1045C : rd_rsp_data <= 32'h00000400;
        16'h10460 : rd_rsp_data <= 32'h00005105;
        16'h107F0 : rd_rsp_data <= 32'h01000208;
        16'h107F4 : rd_rsp_data <= 32'h00000400;
        16'h107F8 : rd_rsp_data <= 32'h0100021A;
        16'h107FC : rd_rsp_data <= 32'h00000400;
        16'h10C00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10C9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10CFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10D9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10DFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10E9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10ECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10ED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10ED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10ED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10EFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10F9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h10FFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11000 : rd_rsp_data <= 32'h01000208;
        16'h11004 : rd_rsp_data <= 32'h00000400;
        16'h11008 : rd_rsp_data <= 32'h0100021A;
        16'h1100C : rd_rsp_data <= 32'h00000400;
        16'h11010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11018 : rd_rsp_data <= 32'h01000208;
        16'h1101C : rd_rsp_data <= 32'h00000400;
        16'h11020 : rd_rsp_data <= 32'h0100020A;
        16'h11024 : rd_rsp_data <= 32'h00000400;
        16'h11028 : rd_rsp_data <= 32'h0100020A;
        16'h1102C : rd_rsp_data <= 32'h00000400;
        16'h11030 : rd_rsp_data <= 32'h01000208;
        16'h11034 : rd_rsp_data <= 32'h00000400;
        16'h11038 : rd_rsp_data <= 32'h0100021B;
        16'h1103C : rd_rsp_data <= 32'h00000400;
        16'h11040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11048 : rd_rsp_data <= 32'h00080008;
        16'h1104C : rd_rsp_data <= 32'h00040001;
        16'h11050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1105C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11068 : rd_rsp_data <= 32'h00000A10;
        16'h1106C : rd_rsp_data <= 32'h00100100;
        16'h11070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11078 : rd_rsp_data <= 32'h000003C0;
        16'h1107C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11080 : rd_rsp_data <= 32'h07040303;
        16'h11084 : rd_rsp_data <= 32'h00000303;
        16'h11088 : rd_rsp_data <= 32'h00000303;
        16'h1108C : rd_rsp_data <= 32'h00000303;
        16'h11090 : rd_rsp_data <= 32'h00000704;
        16'h11098 : rd_rsp_data <= 32'h08040303;
        16'h1109C : rd_rsp_data <= 32'h08040303;
        16'h110A0 : rd_rsp_data <= 32'h00000303;
        16'h110A4 : rd_rsp_data <= 32'h00000303;
        16'h110A8 : rd_rsp_data <= 32'h00001008;
        16'h110B0 : rd_rsp_data <= 32'h05030303;
        16'h110B4 : rd_rsp_data <= 32'h00000303;
        16'h110B8 : rd_rsp_data <= 32'h00000303;
        16'h110BC : rd_rsp_data <= 32'h00000303;
        16'h110C0 : rd_rsp_data <= 32'h00000503;
        16'h110C8 : rd_rsp_data <= 32'h05050303;
        16'h110CC : rd_rsp_data <= 32'h00000303;
        16'h110D0 : rd_rsp_data <= 32'h00000303;
        16'h110D4 : rd_rsp_data <= 32'h00000303;
        16'h110D8 : rd_rsp_data <= 32'h00000505;
        16'h110E0 : rd_rsp_data <= 32'h08080303;
        16'h110E4 : rd_rsp_data <= 32'h08080303;
        16'h110E8 : rd_rsp_data <= 32'h00000303;
        16'h110EC : rd_rsp_data <= 32'h00000303;
        16'h110F0 : rd_rsp_data <= 32'h00011010;
        16'h11100 : rd_rsp_data <= 32'h0002FD32;
        16'h11120 : rd_rsp_data <= 32'h00003910;
        16'h11140 : rd_rsp_data <= 32'h22D1C19B;
        16'h11160 : rd_rsp_data <= 32'h1867FC49;
        16'h11180 : rd_rsp_data <= 32'h00002828;
        16'h11184 : rd_rsp_data <= 32'h0000FF00;
        16'h11450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11800 : rd_rsp_data <= 32'h01000208;
        16'h11804 : rd_rsp_data <= 32'h00000400;
        16'h11808 : rd_rsp_data <= 32'h0100021A;
        16'h1180C : rd_rsp_data <= 32'h00000400;
        16'h11810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11818 : rd_rsp_data <= 32'h01000208;
        16'h1181C : rd_rsp_data <= 32'h00000400;
        16'h11820 : rd_rsp_data <= 32'h0100020A;
        16'h11824 : rd_rsp_data <= 32'h00000400;
        16'h11828 : rd_rsp_data <= 32'h0100020A;
        16'h1182C : rd_rsp_data <= 32'h00000400;
        16'h11830 : rd_rsp_data <= 32'h01000208;
        16'h11834 : rd_rsp_data <= 32'h00000400;
        16'h11838 : rd_rsp_data <= 32'h0100021B;
        16'h1183C : rd_rsp_data <= 32'h00000400;
        16'h11840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11848 : rd_rsp_data <= 32'h00080008;
        16'h1184C : rd_rsp_data <= 32'h00040001;
        16'h11850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1185C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11868 : rd_rsp_data <= 32'h00000A10;
        16'h1186C : rd_rsp_data <= 32'h00100100;
        16'h11870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11878 : rd_rsp_data <= 32'h000003C0;
        16'h1187C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11880 : rd_rsp_data <= 32'h07040303;
        16'h11884 : rd_rsp_data <= 32'h00000303;
        16'h11888 : rd_rsp_data <= 32'h00000303;
        16'h1188C : rd_rsp_data <= 32'h00000303;
        16'h11890 : rd_rsp_data <= 32'h00000704;
        16'h11898 : rd_rsp_data <= 32'h08040303;
        16'h1189C : rd_rsp_data <= 32'h08040303;
        16'h118A0 : rd_rsp_data <= 32'h00000303;
        16'h118A4 : rd_rsp_data <= 32'h00000303;
        16'h118A8 : rd_rsp_data <= 32'h00001008;
        16'h118B0 : rd_rsp_data <= 32'h05030303;
        16'h118B4 : rd_rsp_data <= 32'h00000303;
        16'h118B8 : rd_rsp_data <= 32'h00000303;
        16'h118BC : rd_rsp_data <= 32'h00000303;
        16'h118C0 : rd_rsp_data <= 32'h00000503;
        16'h118C8 : rd_rsp_data <= 32'h05050303;
        16'h118CC : rd_rsp_data <= 32'h00000303;
        16'h118D0 : rd_rsp_data <= 32'h00000303;
        16'h118D4 : rd_rsp_data <= 32'h00000303;
        16'h118D8 : rd_rsp_data <= 32'h00000505;
        16'h118E0 : rd_rsp_data <= 32'h08080303;
        16'h118E4 : rd_rsp_data <= 32'h08080303;
        16'h118E8 : rd_rsp_data <= 32'h00000303;
        16'h118EC : rd_rsp_data <= 32'h00000303;
        16'h118F0 : rd_rsp_data <= 32'h00011010;
        16'h11900 : rd_rsp_data <= 32'h0002FD2D;
        16'h11920 : rd_rsp_data <= 32'h00003916;
        16'h11940 : rd_rsp_data <= 32'h24C32C0F;
        16'h11960 : rd_rsp_data <= 32'h18BA9413;
        16'h11980 : rd_rsp_data <= 32'h00002828;
        16'h11984 : rd_rsp_data <= 32'h0000FF00;
        16'h11C50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h11C54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12000 : rd_rsp_data <= 32'h01000208;
        16'h12004 : rd_rsp_data <= 32'h00000400;
        16'h12008 : rd_rsp_data <= 32'h0100021A;
        16'h1200C : rd_rsp_data <= 32'h00000400;
        16'h12010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12018 : rd_rsp_data <= 32'h01000208;
        16'h1201C : rd_rsp_data <= 32'h00000400;
        16'h12020 : rd_rsp_data <= 32'h0100020A;
        16'h12024 : rd_rsp_data <= 32'h00000400;
        16'h12028 : rd_rsp_data <= 32'h0100020A;
        16'h1202C : rd_rsp_data <= 32'h00000400;
        16'h12030 : rd_rsp_data <= 32'h01000208;
        16'h12034 : rd_rsp_data <= 32'h00000400;
        16'h12038 : rd_rsp_data <= 32'h0100020A;
        16'h1203C : rd_rsp_data <= 32'h00000400;
        16'h12040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12048 : rd_rsp_data <= 32'h01000208;
        16'h1204C : rd_rsp_data <= 32'h00000400;
        16'h12050 : rd_rsp_data <= 32'h0100021B;
        16'h12054 : rd_rsp_data <= 32'h00000400;
        16'h12058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1205C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12060 : rd_rsp_data <= 32'h00080008;
        16'h12064 : rd_rsp_data <= 32'h00040001;
        16'h12068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1206C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12080 : rd_rsp_data <= 32'h00000A10;
        16'h12084 : rd_rsp_data <= 32'h00100100;
        16'h12088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1208C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12090 : rd_rsp_data <= 32'h000003C0;
        16'h12094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12098 : rd_rsp_data <= 32'h09050303;
        16'h1209C : rd_rsp_data <= 32'h09050303;
        16'h120A0 : rd_rsp_data <= 32'h00000303;
        16'h120A4 : rd_rsp_data <= 32'h00000303;
        16'h120A8 : rd_rsp_data <= 32'h0000120A;
        16'h120B0 : rd_rsp_data <= 32'h09050303;
        16'h120B4 : rd_rsp_data <= 32'h09050303;
        16'h120B8 : rd_rsp_data <= 32'h00000303;
        16'h120BC : rd_rsp_data <= 32'h00000303;
        16'h120C0 : rd_rsp_data <= 32'h0000120A;
        16'h120C8 : rd_rsp_data <= 32'h0A050303;
        16'h120CC : rd_rsp_data <= 32'h00000303;
        16'h120D0 : rd_rsp_data <= 32'h00000303;
        16'h120D4 : rd_rsp_data <= 32'h0A080303;
        16'h120D8 : rd_rsp_data <= 32'h0000140D;
        16'h120E0 : rd_rsp_data <= 32'h0A050303;
        16'h120E4 : rd_rsp_data <= 32'h00000303;
        16'h120E8 : rd_rsp_data <= 32'h00000303;
        16'h120EC : rd_rsp_data <= 32'h0A080303;
        16'h120F0 : rd_rsp_data <= 32'h0000140D;
        16'h120F8 : rd_rsp_data <= 32'h00000303;
        16'h120FC : rd_rsp_data <= 32'h00000303;
        16'h12100 : rd_rsp_data <= 32'h00000303;
        16'h12104 : rd_rsp_data <= 32'h05040303;
        16'h12108 : rd_rsp_data <= 32'h00010405;
        16'h12110 : rd_rsp_data <= 32'h00000303;
        16'h12114 : rd_rsp_data <= 32'h00000303;
        16'h12118 : rd_rsp_data <= 32'h00000303;
        16'h1211C : rd_rsp_data <= 32'h05040303;
        16'h12120 : rd_rsp_data <= 32'h00010405;
        16'h12128 : rd_rsp_data <= 32'h0F0E0303;
        16'h1212C : rd_rsp_data <= 32'h0F0E0303;
        16'h12130 : rd_rsp_data <= 32'h00000303;
        16'h12134 : rd_rsp_data <= 32'h00000303;
        16'h12138 : rd_rsp_data <= 32'h00011C1E;
        16'h12140 : rd_rsp_data <= 32'h0F0E0303;
        16'h12144 : rd_rsp_data <= 32'h0F0E0303;
        16'h12148 : rd_rsp_data <= 32'h00000303;
        16'h1214C : rd_rsp_data <= 32'h00000303;
        16'h12150 : rd_rsp_data <= 32'h00011C1E;
        16'h12158 : rd_rsp_data <= 32'h00010000;
        16'h1215C : rd_rsp_data <= 32'h52800000;
        16'h12160 : rd_rsp_data <= 32'h03082404;
        16'h1216C : rd_rsp_data <= 32'h00000004;
        16'h12170 : rd_rsp_data <= 32'hAD7FFFFF;
        16'h12174 : rd_rsp_data <= 32'h00000004;
        16'h12178 : rd_rsp_data <= 32'h00000001;
        16'h12198 : rd_rsp_data <= 32'h0002FD32;
        16'h121B8 : rd_rsp_data <= 32'h00003910;
        16'h121D8 : rd_rsp_data <= 32'h0002FD2D;
        16'h121F8 : rd_rsp_data <= 32'h00003916;
        16'h12200 : rd_rsp_data <= 32'h367E5906;
        16'h12204 : rd_rsp_data <= 32'h0000000F;
        16'h12220 : rd_rsp_data <= 32'h4CE4FFC7;
        16'h12224 : rd_rsp_data <= 32'h00000003;
        16'h12240 : rd_rsp_data <= 32'h39EFB4C3;
        16'h12244 : rd_rsp_data <= 32'h0000000F;
        16'h12260 : rd_rsp_data <= 32'h4D5C0928;
        16'h12264 : rd_rsp_data <= 32'h00000003;
        16'h12280 : rd_rsp_data <= 32'h00002828;
        16'h12284 : rd_rsp_data <= 32'h0000FF00;
        16'h12468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1246C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1280C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1281C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1282C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1283C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1284C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1285C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1286C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1287C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1288C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1289C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h128FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1290C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1291C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1292C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1293C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1294C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1295C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1296C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1297C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1298C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1299C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h129FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12A9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12ABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12ACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12ADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12AFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12B9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12BFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12C9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12CFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12D9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12DFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12E9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12ECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12ED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12ED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12ED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12EFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12F9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h12FFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1300C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1301C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1302C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1303C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1304C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1305C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1306C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1307C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1308C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1309C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h130FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1310C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1311C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1312C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1313C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1314C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1315C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1316C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1317C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1318C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1319C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h131FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1320C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1321C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1322C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1323C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1324C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1325C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1326C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1327C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1328C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1329C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h132FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1330C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1331C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1332C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1333C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1334C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1335C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1336C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1337C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1338C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1339C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h133FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1340C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1341C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1342C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1343C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1344C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1345C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1346C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1347C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1348C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1349C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h134FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1350C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1351C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1352C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1353C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1354C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1355C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1356C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1357C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1358C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1359C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h135FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1360C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1361C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1362C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1363C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1364C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1365C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1366C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1367C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1368C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1369C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h136FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1370C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1371C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1372C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1373C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1374C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1375C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1376C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1377C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1378C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1379C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h137FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1380C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1381C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1382C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1383C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1384C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1385C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1386C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1387C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1388C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1389C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h138FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1390C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1391C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1392C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1393C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1394C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1395C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1396C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1397C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1398C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1399C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h139FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13A9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13ABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13ACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13ADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13AFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13B9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13BFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13C9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13CFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13D9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13DFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13E9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13ECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13ED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13ED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13ED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13EFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13F9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h13FFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1400C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1401C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1402C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1403C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1404C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1405C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1406C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1407C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1408C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1409C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h140FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1410C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1411C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1412C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1413C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1414C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1415C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1416C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1417C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1418C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1419C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h141FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1420C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1421C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1422C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1423C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1424C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1425C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1426C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1427C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1428C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1429C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h142FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1430C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1431C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1432C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1433C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1434C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1435C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1436C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1437C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1438C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1439C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h143FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1440C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1441C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1442C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1443C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1444C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1445C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1446C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1447C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1448C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1449C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h144FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1450C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1451C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1452C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1453C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1454C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1455C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1456C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1457C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1458C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1459C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h145FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1460C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1461C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1462C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1463C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1464C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1465C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1466C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1467C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1468C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1469C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h146FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1470C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1471C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1472C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1473C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1474C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1475C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1476C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1477C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1478C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1479C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h147FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1480C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1481C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1482C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1483C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1484C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1485C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1486C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1487C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1488C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1489C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h148FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1490C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1491C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1492C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1493C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1494C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1495C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1496C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1497C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1498C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1499C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h149FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14A9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14ABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14ACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14ADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14AFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14B9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14BFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14C9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14CFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14D9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14DFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14E9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14ECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14ED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14ED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14ED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14EFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14F9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h14FFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1500C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1501C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1502C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1503C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1504C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1505C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1506C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1507C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1508C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1509C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h150FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1510C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1511C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1512C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1513C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1514C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1515C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1516C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1517C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1518C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1519C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h151FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1520C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1521C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1522C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1523C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1524C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1525C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1526C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1527C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1528C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1529C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h152FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1530C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1531C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1532C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1533C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1534C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1535C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1536C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1537C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1538C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1539C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h153FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1540C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1541C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1542C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1543C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1544C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1545C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1546C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1547C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1548C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1549C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h154FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1550C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1551C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1552C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1553C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1554C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1555C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1556C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1557C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1558C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1559C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h155FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1560C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1561C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1562C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1563C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1564C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1565C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1566C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1567C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1568C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1569C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h156FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1570C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1571C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1572C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1573C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1574C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1575C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1576C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1577C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1578C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1579C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h157FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1580C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1581C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1582C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1583C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1584C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1585C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1586C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1587C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1588C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1589C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h158FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1590C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1591C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1592C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1593C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1594C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1595C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1596C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1597C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1598C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1599C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h159FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15A9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15ABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15ACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15ADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15AFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15B9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15BFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15C9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15CFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15D9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15DFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15E9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15ECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15ED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15ED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15ED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15EFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15F9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h15FFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1600C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1601C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1602C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1603C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1604C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1605C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1606C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1607C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1608C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1609C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h160FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1610C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1611C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1612C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1613C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1614C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1615C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1616C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1617C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1618C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1619C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h161FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1620C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1621C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1622C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1623C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1624C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1625C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1626C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1627C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1628C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1629C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h162FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1630C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1631C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1632C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1633C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1634C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1635C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1636C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1637C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1638C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1639C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h163FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1640C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1641C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1642C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1643C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1644C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1645C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1646C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1647C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1648C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1649C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h164FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1650C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1651C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1652C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1653C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1654C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1655C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1656C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1657C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1658C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1659C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h165FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1660C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1661C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1662C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1663C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1664C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1665C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1666C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1667C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1668C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1669C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h166FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1670C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1671C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1672C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1673C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1674C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1675C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1676C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1677C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1678C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1679C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h167FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1680C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1681C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1682C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1683C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1684C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1685C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1686C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1687C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1688C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1689C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h168FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1690C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1691C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1692C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1693C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1694C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1695C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1696C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1697C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1698C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1699C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h169FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16A9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16ABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16ACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16ADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16AFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16B9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16BFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16C9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16CFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16D9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16DFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16E9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16ECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16ED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16ED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16ED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16EFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16F9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h16FFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1700C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1701C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1702C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1703C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1704C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1705C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1706C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1707C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1708C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1709C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h170FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1710C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1711C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1712C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1713C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1714C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1715C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1716C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1717C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1718C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1719C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h171FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1720C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1721C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1722C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1723C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1724C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1725C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1726C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1727C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1728C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1729C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h172FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1730C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1731C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1732C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1733C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1734C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1735C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1736C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1737C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1738C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1739C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h173FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1740C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1741C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1742C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1743C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1744C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1745C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1746C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1747C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1748C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1749C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h174FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1750C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1751C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1752C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1753C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1754C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1755C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1756C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1757C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1758C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1759C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h175FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1760C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1761C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1762C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1763C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1764C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1765C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1766C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1767C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1768C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1769C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h176FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1770C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1771C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1772C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1773C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1774C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1775C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1776C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1777C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1778C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1779C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h177FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1780C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1781C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1782C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1783C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1784C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1785C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1786C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1787C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1788C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1789C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h178FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1790C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1791C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1792C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1793C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1794C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1795C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1796C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1797C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1798C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1799C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h179FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17A9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17ABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17ACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17ADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17AFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17B9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17BFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17C9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17CFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17D9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17DFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17E9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17ECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17ED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17ED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17ED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17EFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17F9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h17FFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1800C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1801C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1802C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1803C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1804C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1805C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1806C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1807C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1808C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1809C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h180FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1810C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1811C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1812C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1813C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1814C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1815C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1816C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1817C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1818C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1819C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h181FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1820C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1821C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1822C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1823C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1824C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1825C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1826C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1827C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1828C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1829C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h182FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1830C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1831C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1832C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1833C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1834C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1835C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1836C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1837C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1838C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1839C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h183FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1840C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1841C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1842C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1843C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1844C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1845C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1846C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1847C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1848C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1849C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h184FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1850C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1851C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1852C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1853C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1854C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1855C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1856C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1857C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1858C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1859C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h185FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1860C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1861C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1862C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1863C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1864C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1865C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1866C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1867C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1868C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1869C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h186FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1870C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1871C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1872C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1873C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1874C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1875C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1876C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1877C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1878C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1879C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h187FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1880C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1881C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1882C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1883C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1884C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1885C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1886C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1887C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1888C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1889C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h188FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1890C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1891C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1892C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1893C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1894C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1895C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1896C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1897C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1898C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1899C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h189FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18A9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18ABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18ACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18ADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18AFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18B9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18BFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18C9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18CFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18D9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18DFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18E9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18ECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18ED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18ED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18ED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18EFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18F9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h18FFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1900C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1901C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1902C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1903C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1904C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1905C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1906C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1907C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1908C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1909C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h190FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1910C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1911C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1912C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1913C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1914C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1915C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1916C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1917C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1918C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1919C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h191FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1920C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1921C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1922C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1923C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1924C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1925C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1926C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1927C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1928C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1929C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h192FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1930C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1931C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1932C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1933C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1934C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1935C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1936C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1937C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1938C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1939C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h193FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1940C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1941C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1942C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1943C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1944C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1945C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1946C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1947C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1948C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1949C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h194FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1950C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1951C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1952C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1953C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1954C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1955C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1956C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1957C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1958C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1959C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h195FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1960C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1961C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1962C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1963C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1964C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1965C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1966C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1967C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1968C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1969C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h196FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1970C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1971C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1972C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1973C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1974C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1975C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1976C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1977C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1978C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1979C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h197FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1980C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1981C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1982C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1983C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1984C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1985C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1986C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1987C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1988C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1989C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h198FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1990C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1991C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1992C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1993C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1994C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1995C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1996C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1997C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1998C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1999C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h199FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19A9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19ABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19ACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19ADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19AFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19B9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19BFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19C9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19CFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19D9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19DFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19E9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19ECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19ED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19ED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19ED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19EFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19F9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h19FFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A00C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A01C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A02C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A03C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A04C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A05C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A06C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A07C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A08C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A09C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A0FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A10C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A11C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A12C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A13C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A14C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A15C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A16C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A17C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A18C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A19C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A1FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A20C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A21C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A22C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A23C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A24C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A25C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A26C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A27C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A28C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A29C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A2FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A30C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A31C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A32C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A33C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A34C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A35C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A36C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A37C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A38C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A39C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A3FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A40C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A41C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A42C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A43C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A44C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A45C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A46C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A47C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A48C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A49C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A4FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A50C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A51C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A52C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A53C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A54C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A55C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A56C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A57C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A58C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A59C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A5FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A60C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A61C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A62C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A63C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A64C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A65C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A66C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A67C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A68C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A69C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A6FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A70C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A71C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A72C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A73C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A74C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A75C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A76C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A77C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A78C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A79C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A7FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A80C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A81C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A82C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A83C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A84C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A85C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A86C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A87C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A88C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A89C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A8FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A90C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A91C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A92C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A93C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A94C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A95C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A96C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A97C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A98C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A99C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1A9FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AA9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AAFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AB9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ABFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AC9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ACFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AD9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1ADFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AE9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AEFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AF9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1AFFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B00C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B01C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B02C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B03C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B04C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B05C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B06C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B07C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B08C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B09C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B0FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B10C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B11C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B12C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B13C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B14C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B15C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B16C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B17C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B18C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B19C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B1FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B20C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B21C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B22C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B23C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B24C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B25C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B26C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B27C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B28C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B29C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B2FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B30C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B31C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B32C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B33C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B34C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B35C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B36C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B37C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B38C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B39C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B3FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B40C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B41C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B42C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B43C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B44C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B45C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B46C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B47C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B48C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B49C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B4FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B50C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B51C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B52C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B53C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B54C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B55C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B56C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B57C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B58C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B59C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B5FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B60C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B61C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B62C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B63C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B64C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B65C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B66C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B67C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B68C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B69C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B6FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B70C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B71C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B72C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B73C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B74C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B75C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B76C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B77C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B78C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B79C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B7FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B80C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B81C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B82C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B83C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B84C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B85C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B86C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B87C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B88C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B89C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B8FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B90C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B91C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B92C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B93C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B94C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B95C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B96C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B97C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B98C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B99C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1B9FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BA9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BAFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BB9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BBFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BC9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BCFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BD9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BDFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BE9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BEFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BF9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1BFFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C000 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C004 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C00C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C010 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C014 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C018 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C01C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C020 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C024 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C028 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C02C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C030 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C034 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C038 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C03C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C040 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C044 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C048 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C04C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C050 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C054 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C058 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C05C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C060 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C064 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C068 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C06C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C070 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C074 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C078 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C07C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C080 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C084 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C088 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C08C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C090 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C094 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C098 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C09C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C0FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C100 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C104 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C10C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C110 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C114 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C118 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C11C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C120 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C124 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C128 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C12C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C130 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C134 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C138 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C13C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C140 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C144 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C148 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C14C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C150 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C154 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C158 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C15C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C160 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C164 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C168 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C16C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C170 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C174 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C178 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C17C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C180 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C184 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C188 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C18C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C190 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C194 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C198 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C19C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C1FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C200 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C204 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C20C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C210 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C214 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C218 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C21C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C220 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C224 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C228 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C22C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C230 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C234 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C238 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C23C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C240 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C244 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C248 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C24C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C250 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C254 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C258 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C25C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C260 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C264 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C268 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C26C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C270 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C274 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C278 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C27C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C280 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C284 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C288 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C28C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C290 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C294 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C298 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C29C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C2FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C300 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C304 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C30C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C310 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C314 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C318 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C31C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C320 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C324 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C328 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C32C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C330 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C334 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C338 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C33C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C340 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C344 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C348 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C34C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C350 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C354 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C358 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C35C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C360 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C364 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C368 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C36C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C370 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C374 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C378 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C37C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C380 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C384 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C388 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C38C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C390 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C394 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C398 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C39C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C3FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C40C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C41C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C42C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C43C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C44C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C45C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C46C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C47C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C48C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C49C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C4FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C50C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C51C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C52C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C53C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C54C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C55C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C56C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C57C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C58C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C59C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C5FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C60C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C61C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C62C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C63C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C64C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C65C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C66C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C67C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C68C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C69C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C6FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C70C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C71C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C72C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C73C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C74C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C75C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C76C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C77C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C78C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C79C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C7FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C800 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C804 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C808 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C80C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C810 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C814 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C818 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C81C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C820 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C824 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C828 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C82C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C830 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C834 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C838 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C83C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C840 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C844 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C848 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C84C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C850 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C854 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C858 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C85C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C860 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C864 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C868 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C86C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C870 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C874 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C878 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C87C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C880 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C884 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C888 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C88C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C890 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C894 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C898 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C89C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C8FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C900 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C904 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C908 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C90C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C910 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C914 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C918 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C91C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C920 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C924 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C928 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C92C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C930 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C934 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C938 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C93C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C940 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C944 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C948 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C94C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C950 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C954 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C95C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C960 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C964 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C968 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C96C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C970 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C974 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C978 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C97C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C980 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C984 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C988 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C98C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C990 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C994 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C998 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C99C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1C9FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CA9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CABC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CACC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CADC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CAFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CB9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CBFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CC9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CCFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CD9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CDFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CE9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CECC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CED0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CED4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CED8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CEFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF00 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF04 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF08 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF0C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF10 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF14 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF18 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF1C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF20 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF24 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF28 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF2C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF30 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF34 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF38 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF3C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF40 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF44 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF48 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF4C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF50 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF54 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF58 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF5C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF60 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF64 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF68 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF6C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF70 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF74 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF78 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF7C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF80 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF84 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF88 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF8C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF90 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF94 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF98 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CF9C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFA0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFA4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFA8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFAC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFB0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFB4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFB8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFBC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFC0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFC4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFC8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFCC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFD0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFD4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFD8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFDC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFE0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFE4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFE8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFEC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFF0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFF4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFF8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1CFFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D000 : rd_rsp_data <= 32'h01000208;
        16'h1D004 : rd_rsp_data <= 32'h00000400;
        16'h1D008 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D00C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D010 : rd_rsp_data <= 32'h0100021A;
        16'h1D014 : rd_rsp_data <= 32'h00000400;
        16'h1D01C : rd_rsp_data <= 32'h00001800;
        16'h1D028 : rd_rsp_data <= 32'h01040000;
        16'h1D030 : rd_rsp_data <= 32'h00411421;
        16'h1D038 : rd_rsp_data <= 32'h00010101;
        16'h1D040 : rd_rsp_data <= 32'h0000AA55;
        16'h1D044 : rd_rsp_data <= 32'h0000AA55;
        16'h1D048 : rd_rsp_data <= 32'h0000AA55;
        16'h1D050 : rd_rsp_data <= 32'h01010100;
        16'h1D058 : rd_rsp_data <= 32'h80000000;
        16'h1D05C : rd_rsp_data <= 32'h80000000;
        16'h1D060 : rd_rsp_data <= 32'h80000000;
        16'h1D100 : rd_rsp_data <= 32'h01000208;
        16'h1D104 : rd_rsp_data <= 32'h00000400;
        16'h1D108 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D10C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D110 : rd_rsp_data <= 32'h0100021A;
        16'h1D114 : rd_rsp_data <= 32'h00000400;
        16'h1D11C : rd_rsp_data <= 32'h00001800;
        16'h1D128 : rd_rsp_data <= 32'h00640000;
        16'h1D130 : rd_rsp_data <= 32'h00411421;
        16'h1D138 : rd_rsp_data <= 32'h00010101;
        16'h1D140 : rd_rsp_data <= 32'h0000AA55;
        16'h1D144 : rd_rsp_data <= 32'h0000AA55;
        16'h1D148 : rd_rsp_data <= 32'h0000AA55;
        16'h1D150 : rd_rsp_data <= 32'h01010100;
        16'h1D158 : rd_rsp_data <= 32'h80000000;
        16'h1D15C : rd_rsp_data <= 32'h80000000;
        16'h1D160 : rd_rsp_data <= 32'h80000000;
        16'h1D200 : rd_rsp_data <= 32'h01000208;
        16'h1D204 : rd_rsp_data <= 32'h00000400;
        16'h1D208 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D20C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D210 : rd_rsp_data <= 32'h0100021A;
        16'h1D214 : rd_rsp_data <= 32'h00000400;
        16'h1D21C : rd_rsp_data <= 32'h00001800;
        16'h1D228 : rd_rsp_data <= 32'h01040000;
        16'h1D230 : rd_rsp_data <= 32'h00411421;
        16'h1D238 : rd_rsp_data <= 32'h00010101;
        16'h1D240 : rd_rsp_data <= 32'h0000AA55;
        16'h1D244 : rd_rsp_data <= 32'h0000AA55;
        16'h1D248 : rd_rsp_data <= 32'h0000AA55;
        16'h1D250 : rd_rsp_data <= 32'h01010100;
        16'h1D258 : rd_rsp_data <= 32'h80000000;
        16'h1D25C : rd_rsp_data <= 32'h80000000;
        16'h1D260 : rd_rsp_data <= 32'h80000000;
        16'h1D300 : rd_rsp_data <= 32'h01000208;
        16'h1D304 : rd_rsp_data <= 32'h00000400;
        16'h1D308 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D30C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D310 : rd_rsp_data <= 32'h0100021A;
        16'h1D314 : rd_rsp_data <= 32'h00000400;
        16'h1D31C : rd_rsp_data <= 32'h00001800;
        16'h1D328 : rd_rsp_data <= 32'h00640000;
        16'h1D330 : rd_rsp_data <= 32'h00411421;
        16'h1D338 : rd_rsp_data <= 32'h00010101;
        16'h1D340 : rd_rsp_data <= 32'h0000AA55;
        16'h1D344 : rd_rsp_data <= 32'h0000AA55;
        16'h1D348 : rd_rsp_data <= 32'h0000AA55;
        16'h1D350 : rd_rsp_data <= 32'h01010100;
        16'h1D358 : rd_rsp_data <= 32'h80000000;
        16'h1D35C : rd_rsp_data <= 32'h80000000;
        16'h1D360 : rd_rsp_data <= 32'h80000000;
        16'h1D400 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D404 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D408 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D40C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D410 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D414 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D418 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D41C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D420 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D424 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D428 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D42C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D430 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D434 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D438 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D43C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D440 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D444 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D448 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D44C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D450 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D454 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D458 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D45C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D460 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D464 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D468 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D46C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D470 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D474 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D478 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D47C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D480 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D484 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D488 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D48C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D490 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D494 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D498 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D49C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D4FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D500 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D504 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D508 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D50C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D510 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D514 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D518 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D51C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D520 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D524 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D528 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D52C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D530 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D534 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D538 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D53C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D540 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D544 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D548 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D54C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D550 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D554 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D558 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D55C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D560 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D564 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D568 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D56C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D570 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D574 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D578 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D57C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D580 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D584 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D588 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D58C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D590 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D594 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D598 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D59C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D5FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D600 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D604 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D608 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D60C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D610 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D614 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D618 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D61C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D620 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D624 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D628 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D62C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D630 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D634 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D638 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D63C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D640 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D644 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D648 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D64C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D650 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D654 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D658 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D65C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D660 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D664 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D668 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D66C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D670 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D674 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D678 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D67C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D680 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D684 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D688 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D68C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D690 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D694 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D698 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D69C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D6FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D700 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D704 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D708 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D70C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D710 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D714 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D718 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D71C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D720 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D724 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D728 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D72C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D730 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D734 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D738 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D73C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D740 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D744 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D748 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D74C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D750 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D754 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D758 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D75C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D760 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D764 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D768 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D76C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D770 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D774 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D778 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D77C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D780 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D784 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D788 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D78C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D790 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D794 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D798 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D79C : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7A0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7A4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7A8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7AC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7B0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7B4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7B8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7BC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7C0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7C4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7C8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7CC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7D0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7D4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7D8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7DC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7E0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7E4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7E8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7EC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7F0 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7F4 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7F8 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D7FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D800 : rd_rsp_data <= 32'h08008001;
        16'h1D804 : rd_rsp_data <= 32'h00000100;
        16'h1D808 : rd_rsp_data <= 32'h00000100;
        16'h1D80C : rd_rsp_data <= 32'hD0000088;
        16'h1D810 : rd_rsp_data <= 32'hD0000088;
        16'h1D814 : rd_rsp_data <= 32'h00000002;
        16'h1D81C : rd_rsp_data <= 32'h00018200;
        16'h1D824 : rd_rsp_data <= 32'h130C3200;
        16'h1D830 : rd_rsp_data <= 32'h004000AA;
        16'h1D83C : rd_rsp_data <= 32'h00010820;
        16'h1D840 : rd_rsp_data <= 32'h874C3B28;
        16'h1D844 : rd_rsp_data <= 32'h00000012;
        16'h1D858 : rd_rsp_data <= 32'h3C46E0BA;
        16'h1D85C : rd_rsp_data <= 32'h0000000F;
        16'h1D860 : rd_rsp_data <= 32'h00010200;
        16'h1D874 : rd_rsp_data <= 32'h00000010;
        16'h1D878 : rd_rsp_data <= 32'h00001844;
        16'h1D87C : rd_rsp_data <= 32'h00001844;
        16'h1D880 : rd_rsp_data <= 32'h24504030;
        16'h1D890 : rd_rsp_data <= 32'hFFF00000;
        16'h1D894 : rd_rsp_data <= 32'h0000007F;
        16'h1D8A0 : rd_rsp_data <= 32'h488EDDE0;
        16'h1D8A4 : rd_rsp_data <= 32'h00000003;
        16'h1D8A8 : rd_rsp_data <= 32'hFDDE557B;
        16'h1D8AC : rd_rsp_data <= 32'h00000023;
        16'h1D8BC : rd_rsp_data <= 32'h00100000;
        16'h1D930 : rd_rsp_data <= 32'h70B40384;
        16'h1D934 : rd_rsp_data <= 32'h0400B05A;
        16'h1D938 : rd_rsp_data <= 32'h0000000F;
        16'h1D93C : rd_rsp_data <= 32'h00301C1C;
        16'h1D954 : rd_rsp_data <= 32'h00300100;
        16'h1D958 : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1D95C : rd_rsp_data <= 32'h00000001;
        16'h1D960 : rd_rsp_data <= 32'h038400E1;
        16'h1D964 : rd_rsp_data <= 32'h0000005A;
        16'h1D968 : rd_rsp_data <= 32'h0001407D;
        16'h1D96C : rd_rsp_data <= 32'h00000001;
        16'h1D974 : rd_rsp_data <= 32'h000000C6;
        16'h1D9B4 : rd_rsp_data <= 32'h0000001F;
        16'h1D9B8 : rd_rsp_data <= 32'h00000107;
        16'h1E000 : rd_rsp_data <= 32'h27422027;
        16'h1E004 : rd_rsp_data <= 32'h01393075;
        16'h1E008 : rd_rsp_data <= 32'h49041828;
        16'h1E00C : rd_rsp_data <= 32'h0E0E088C;
        16'h1E010 : rd_rsp_data <= 32'h16141212;
        16'h1E014 : rd_rsp_data <= 32'h18306C48;
        16'h1E018 : rd_rsp_data <= 32'h0E0E081A;
        16'h1E01C : rd_rsp_data <= 32'h003FF020;
        16'h1E020 : rd_rsp_data <= 32'h19191944;
        16'h1E024 : rd_rsp_data <= 32'h19191919;
        16'h1E028 : rd_rsp_data <= 32'h80000020;
        16'h1E02C : rd_rsp_data <= 32'h4E000200;
        16'h1E034 : rd_rsp_data <= 32'h060101A8;
        16'h1E038 : rd_rsp_data <= 32'h00000C00;
        16'h1E040 : rd_rsp_data <= 32'h000201A8;
        16'h1E044 : rd_rsp_data <= 32'h00000200;
        16'h1E050 : rd_rsp_data <= 32'h060E8912;
        16'h1E054 : rd_rsp_data <= 32'h12068076;
        16'h1E068 : rd_rsp_data <= 32'h103B2838;
        16'h1E06C : rd_rsp_data <= 32'h16404030;
        16'h1E070 : rd_rsp_data <= 32'h26280000;
        16'h1E074 : rd_rsp_data <= 32'h00000080;
        16'h1E078 : rd_rsp_data <= 32'h00300004;
        16'h1E088 : rd_rsp_data <= 32'h8FC00029;
        16'h1E08C : rd_rsp_data <= 32'h0C008484;
        16'h1E090 : rd_rsp_data <= 32'h0C180810;
        16'h1E094 : rd_rsp_data <= 32'h08100408;
        16'h1E098 : rd_rsp_data <= 32'h040C0206;
        16'h1E0A0 : rd_rsp_data <= 32'hD4CA450A;
        16'h1E0A8 : rd_rsp_data <= 32'h02540040;
        16'h1E0AC : rd_rsp_data <= 32'h0281284B;
        16'h1E0B0 : rd_rsp_data <= 32'h0000000F;
        16'h1E0B8 : rd_rsp_data <= 32'h08104426;
        16'h1E0C0 : rd_rsp_data <= 32'h00200086;
        16'h1E0C4 : rd_rsp_data <= 32'h800308E2;
        16'h1E0C8 : rd_rsp_data <= 32'h1C483616;
        16'h1E0D0 : rd_rsp_data <= 32'h0000000F;
        16'h1E0D4 : rd_rsp_data <= 32'h0E64E893;
        16'h1E100 : rd_rsp_data <= 32'h80202028;
        16'h1E110 : rd_rsp_data <= 32'h00000056;
        16'h1E114 : rd_rsp_data <= 32'h00020611;
        16'h1E118 : rd_rsp_data <= 32'hFFF080AE;
        16'h1E11C : rd_rsp_data <= 32'h0001B20A;
        16'h1E120 : rd_rsp_data <= 32'h000000E0;
        16'h1E124 : rd_rsp_data <= 32'h00004000;
        16'h1E128 : rd_rsp_data <= 32'h20000000;
        16'h1E12C : rd_rsp_data <= 32'h00000007;
        16'h1E200 : rd_rsp_data <= 32'h30200884;
        16'h1E204 : rd_rsp_data <= 32'h4F3F2F40;
        16'h1E208 : rd_rsp_data <= 32'h5E56B733;
        16'h1E20C : rd_rsp_data <= 32'h00129024;
        16'h1E210 : rd_rsp_data <= 32'h00040844;
        16'h1E214 : rd_rsp_data <= 32'h80C3C3E8;
        16'h1E218 : rd_rsp_data <= 32'h1B000036;
        16'h1E21C : rd_rsp_data <= 32'h3F001B1B;
        16'h1E220 : rd_rsp_data <= 32'h33333939;
        16'h1E224 : rd_rsp_data <= 32'h0000007F;
        16'h1E3E0 : rd_rsp_data <= 32'h013E9828;
        16'h1E3E4 : rd_rsp_data <= 32'h0000508D;
        16'h1E3F0 : rd_rsp_data <= 32'h01DF23FF;
        16'h1E3F4 : rd_rsp_data <= 32'hB8EF2DCE;
        16'h1E400 : rd_rsp_data <= 32'h11002EC3;
        16'h1E404 : rd_rsp_data <= 32'h0000000F;
        16'h1E40C : rd_rsp_data <= 32'h00000137;
        16'h1E410 : rd_rsp_data <= 32'h00200D05;
        16'h1E418 : rd_rsp_data <= 32'h02020202;
        16'h1E424 : rd_rsp_data <= 32'h00000001;
        16'h1E428 : rd_rsp_data <= 32'h01010101;
        16'h1E42C : rd_rsp_data <= 32'h00101020;
        16'h1E430 : rd_rsp_data <= 32'h23444688;
        16'h1E434 : rd_rsp_data <= 32'h00000008;
        16'h1E438 : rd_rsp_data <= 32'h275A7640;
        16'h1E43C : rd_rsp_data <= 32'h05FC11C5;
        16'h1E440 : rd_rsp_data <= 32'h28000600;
        16'h1E444 : rd_rsp_data <= 32'h00004000;
        16'h1E448 : rd_rsp_data <= 32'h00013880;
        16'h1E44C : rd_rsp_data <= 32'h000004B3;
        16'h1E450 : rd_rsp_data <= 32'h00000012;
        16'h1E454 : rd_rsp_data <= 32'h00000001;
        16'h1E458 : rd_rsp_data <= 32'h00001C00;
        16'h1E46C : rd_rsp_data <= 32'h00000101;
        16'h1E470 : rd_rsp_data <= 32'h00000101;
        16'h1E474 : rd_rsp_data <= 32'h00300E08;
        16'h1E478 : rd_rsp_data <= 32'h00000003;
        16'h1E480 : rd_rsp_data <= 32'h23444688;
        16'h1E484 : rd_rsp_data <= 32'h00000009;
        16'h1E488 : rd_rsp_data <= 32'h0AC4DC14;
        16'h1E494 : rd_rsp_data <= 32'h11311022;
        16'h1E498 : rd_rsp_data <= 32'h23444688;
        16'h1E49C : rd_rsp_data <= 32'h00000008;
        16'h1E4B0 : rd_rsp_data <= 32'h0DC910CB;
        16'h1E4B8 : rd_rsp_data <= 32'h23444688;
        16'h1E4BC : rd_rsp_data <= 32'h0000001B;
        16'h1E4C0 : rd_rsp_data <= 32'h000002C2;
        16'h1E4C4 : rd_rsp_data <= 32'h02000140;
        16'h1E4C8 : rd_rsp_data <= 32'h0C078000;
        16'h1E4D8 : rd_rsp_data <= 32'h854653C3;
        16'h1E4DC : rd_rsp_data <= 32'h56ABF65C;
        16'h1E4FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1E5CC : rd_rsp_data <= 32'h3F000000;
        16'h1E5D0 : rd_rsp_data <= 32'hE0400000;
        16'h1E5D4 : rd_rsp_data <= 32'h26000400;
        16'h1E5E0 : rd_rsp_data <= 32'h00002003;
        16'h1E5E4 : rd_rsp_data <= 32'h0000000F;
        16'h1E5FC : rd_rsp_data <= 32'h08041000;
        16'h1E600 : rd_rsp_data <= 32'h80400000;
        16'h1E604 : rd_rsp_data <= 32'h8040010E;
        16'h1E608 : rd_rsp_data <= 32'h80400201;
        16'h1E60C : rd_rsp_data <= 32'h80400302;
        16'h1E610 : rd_rsp_data <= 32'h80400405;
        16'h1E614 : rd_rsp_data <= 32'h80400503;
        16'h1E618 : rd_rsp_data <= 32'h80400604;
        16'h1E61C : rd_rsp_data <= 32'h80400707;
        16'h1E620 : rd_rsp_data <= 32'h8480080B;
        16'h1E624 : rd_rsp_data <= 32'h8480090C;
        16'h1E628 : rd_rsp_data <= 32'h80400A06;
        16'h1E62C : rd_rsp_data <= 32'h80400B08;
        16'h1E630 : rd_rsp_data <= 32'h80000C00;
        16'h1E634 : rd_rsp_data <= 32'h80000D02;
        16'h1E638 : rd_rsp_data <= 32'h80000E04;
        16'h1E63C : rd_rsp_data <= 32'h80000F05;
        16'h1E640 : rd_rsp_data <= 32'h80001006;
        16'h1E644 : rd_rsp_data <= 32'h80001108;
        16'h1E648 : rd_rsp_data <= 32'h8000120D;
        16'h1E64C : rd_rsp_data <= 32'h8000130E;
        16'h1E650 : rd_rsp_data <= 32'h80001481;
        16'h1E654 : rd_rsp_data <= 32'h80001582;
        16'h1E658 : rd_rsp_data <= 32'h80001683;
        16'h1E65C : rd_rsp_data <= 32'h80001784;
        16'h1E660 : rd_rsp_data <= 32'h80001489;
        16'h1E664 : rd_rsp_data <= 32'h8000158A;
        16'h1E668 : rd_rsp_data <= 32'h8000168B;
        16'h1E66C : rd_rsp_data <= 32'h8000178C;
        16'h1E670 : rd_rsp_data <= 32'h80001491;
        16'h1E674 : rd_rsp_data <= 32'h80001592;
        16'h1E678 : rd_rsp_data <= 32'h80001693;
        16'h1E67C : rd_rsp_data <= 32'h80001794;
        16'h1E680 : rd_rsp_data <= 32'h80001499;
        16'h1E684 : rd_rsp_data <= 32'h8000159A;
        16'h1E688 : rd_rsp_data <= 32'h8000169B;
        16'h1E68C : rd_rsp_data <= 32'h8000179C;
        16'h1E690 : rd_rsp_data <= 32'h800014A1;
        16'h1E694 : rd_rsp_data <= 32'h800015A2;
        16'h1E698 : rd_rsp_data <= 32'h800016A3;
        16'h1E69C : rd_rsp_data <= 32'h800017A4;
        16'h1E6A0 : rd_rsp_data <= 32'h800014A9;
        16'h1E6A4 : rd_rsp_data <= 32'h800015AA;
        16'h1E6A8 : rd_rsp_data <= 32'h800016AB;
        16'h1E6AC : rd_rsp_data <= 32'h800017AC;
        16'h1E6B0 : rd_rsp_data <= 32'h800014B1;
        16'h1E6B4 : rd_rsp_data <= 32'h800015B2;
        16'h1E6B8 : rd_rsp_data <= 32'h800016B3;
        16'h1E6BC : rd_rsp_data <= 32'h800017B4;
        16'h1E6C0 : rd_rsp_data <= 32'h800014B9;
        16'h1E6C4 : rd_rsp_data <= 32'h800015BA;
        16'h1E6C8 : rd_rsp_data <= 32'h800016BB;
        16'h1E6CC : rd_rsp_data <= 32'h800017BC;
        16'h1E6D0 : rd_rsp_data <= 32'h800014C1;
        16'h1E6D4 : rd_rsp_data <= 32'h800015C2;
        16'h1E6D8 : rd_rsp_data <= 32'h800016C3;
        16'h1E6DC : rd_rsp_data <= 32'h800017C4;
        16'h1E6E0 : rd_rsp_data <= 32'h800014C9;
        16'h1E6E4 : rd_rsp_data <= 32'h800015CA;
        16'h1E6E8 : rd_rsp_data <= 32'h800016CB;
        16'h1E6EC : rd_rsp_data <= 32'h800017CC;
        16'h1E6F0 : rd_rsp_data <= 32'h800014D1;
        16'h1E6F4 : rd_rsp_data <= 32'h800015D2;
        16'h1E6F8 : rd_rsp_data <= 32'h800016D3;
        16'h1E6FC : rd_rsp_data <= 32'h800017D4;
        16'h1E700 : rd_rsp_data <= 32'h800014D9;
        16'h1E704 : rd_rsp_data <= 32'h800015DA;
        16'h1E708 : rd_rsp_data <= 32'h800016DB;
        16'h1E70C : rd_rsp_data <= 32'h800017DC;
        16'h1E710 : rd_rsp_data <= 32'h800014E1;
        16'h1E714 : rd_rsp_data <= 32'h800015E2;
        16'h1E718 : rd_rsp_data <= 32'h800016E3;
        16'h1E71C : rd_rsp_data <= 32'h800017E4;
        16'h1E720 : rd_rsp_data <= 32'h800014E9;
        16'h1E724 : rd_rsp_data <= 32'h800015EA;
        16'h1E728 : rd_rsp_data <= 32'h800016EB;
        16'h1E72C : rd_rsp_data <= 32'h800017EC;
        16'h1E730 : rd_rsp_data <= 32'h800014F1;
        16'h1E734 : rd_rsp_data <= 32'h800015F2;
        16'h1E738 : rd_rsp_data <= 32'h800016F3;
        16'h1E73C : rd_rsp_data <= 32'h800017F4;
        16'h1E740 : rd_rsp_data <= 32'h800014F9;
        16'h1E744 : rd_rsp_data <= 32'h800015FA;
        16'h1E748 : rd_rsp_data <= 32'h800016FB;
        16'h1E74C : rd_rsp_data <= 32'h830017FC;
        16'h1E750 : rd_rsp_data <= 32'h80001822;
        16'h1E754 : rd_rsp_data <= 32'h80001923;
        16'h1E758 : rd_rsp_data <= 32'h80001A24;
        16'h1E75C : rd_rsp_data <= 32'h80001B25;
        16'h1E760 : rd_rsp_data <= 32'h80001C26;
        16'h1E764 : rd_rsp_data <= 32'h80001D27;
        16'h1E768 : rd_rsp_data <= 32'h80001E28;
        16'h1E76C : rd_rsp_data <= 32'h80001F2D;
        16'h1E770 : rd_rsp_data <= 32'hC800200A;
        16'h1E774 : rd_rsp_data <= 32'hC8002203;
        16'h1E778 : rd_rsp_data <= 32'h8040240F;
        16'h1E800 : rd_rsp_data <= 32'h27422027;
        16'h1E804 : rd_rsp_data <= 32'h01393075;
        16'h1E808 : rd_rsp_data <= 32'h49041828;
        16'h1E80C : rd_rsp_data <= 32'h0E0E088C;
        16'h1E810 : rd_rsp_data <= 32'h16141212;
        16'h1E814 : rd_rsp_data <= 32'h18306C48;
        16'h1E818 : rd_rsp_data <= 32'h0E0E081A;
        16'h1E81C : rd_rsp_data <= 32'h003FF020;
        16'h1E820 : rd_rsp_data <= 32'h1919193F;
        16'h1E824 : rd_rsp_data <= 32'h19191919;
        16'h1E828 : rd_rsp_data <= 32'h80000020;
        16'h1E82C : rd_rsp_data <= 32'h4E000200;
        16'h1E834 : rd_rsp_data <= 32'h06010138;
        16'h1E838 : rd_rsp_data <= 32'h00000C00;
        16'h1E840 : rd_rsp_data <= 32'h00020138;
        16'h1E844 : rd_rsp_data <= 32'h00000200;
        16'h1E850 : rd_rsp_data <= 32'h060E8912;
        16'h1E854 : rd_rsp_data <= 32'h12068076;
        16'h1E868 : rd_rsp_data <= 32'h103B2838;
        16'h1E86C : rd_rsp_data <= 32'h16404030;
        16'h1E870 : rd_rsp_data <= 32'h26280000;
        16'h1E874 : rd_rsp_data <= 32'h00000080;
        16'h1E878 : rd_rsp_data <= 32'h00300004;
        16'h1E888 : rd_rsp_data <= 32'h8FC00029;
        16'h1E88C : rd_rsp_data <= 32'h0C008484;
        16'h1E890 : rd_rsp_data <= 32'h0C180810;
        16'h1E894 : rd_rsp_data <= 32'h08100408;
        16'h1E898 : rd_rsp_data <= 32'h040C0206;
        16'h1E8A0 : rd_rsp_data <= 32'hD4CA450A;
        16'h1E8A8 : rd_rsp_data <= 32'h02540040;
        16'h1E8AC : rd_rsp_data <= 32'h0281284B;
        16'h1E8B0 : rd_rsp_data <= 32'h0000000F;
        16'h1E8B8 : rd_rsp_data <= 32'h08104426;
        16'h1E8C0 : rd_rsp_data <= 32'h00200086;
        16'h1E8C4 : rd_rsp_data <= 32'h800308E2;
        16'h1E8C8 : rd_rsp_data <= 32'h1C483616;
        16'h1E8D0 : rd_rsp_data <= 32'h0000000F;
        16'h1E8D4 : rd_rsp_data <= 32'h0E64E893;
        16'h1E900 : rd_rsp_data <= 32'h80202028;
        16'h1E910 : rd_rsp_data <= 32'h00000056;
        16'h1E914 : rd_rsp_data <= 32'h00020611;
        16'h1E918 : rd_rsp_data <= 32'hFFF080AE;
        16'h1E91C : rd_rsp_data <= 32'h0001B20A;
        16'h1E920 : rd_rsp_data <= 32'h000000E0;
        16'h1E924 : rd_rsp_data <= 32'h00004000;
        16'h1E928 : rd_rsp_data <= 32'h20000000;
        16'h1E92C : rd_rsp_data <= 32'h00000007;
        16'h1EA00 : rd_rsp_data <= 32'h30200884;
        16'h1EA04 : rd_rsp_data <= 32'h4F3F2F40;
        16'h1EA08 : rd_rsp_data <= 32'h5E56B734;
        16'h1EA0C : rd_rsp_data <= 32'h00129024;
        16'h1EA10 : rd_rsp_data <= 32'h00040844;
        16'h1EA14 : rd_rsp_data <= 32'hC2C3C4E1;
        16'h1EA18 : rd_rsp_data <= 32'h1B000036;
        16'h1EA1C : rd_rsp_data <= 32'h3F001B1B;
        16'h1EA20 : rd_rsp_data <= 32'h33333A3A;
        16'h1EA24 : rd_rsp_data <= 32'h0000007F;
        16'h1EBE0 : rd_rsp_data <= 32'h013E9828;
        16'h1EBE4 : rd_rsp_data <= 32'h0000508D;
        16'h1EBF0 : rd_rsp_data <= 32'h12A0AE5C;
        16'h1EBF4 : rd_rsp_data <= 32'hBFB6D9D1;
        16'h1EC00 : rd_rsp_data <= 32'h11002EC3;
        16'h1EC04 : rd_rsp_data <= 32'h0000000F;
        16'h1EC0C : rd_rsp_data <= 32'h00000137;
        16'h1EC10 : rd_rsp_data <= 32'h00200D05;
        16'h1EC18 : rd_rsp_data <= 32'h02020202;
        16'h1EC24 : rd_rsp_data <= 32'h00000001;
        16'h1EC28 : rd_rsp_data <= 32'h01010101;
        16'h1EC2C : rd_rsp_data <= 32'h00101020;
        16'h1EC30 : rd_rsp_data <= 32'h23444688;
        16'h1EC34 : rd_rsp_data <= 32'h00000008;
        16'h1EC38 : rd_rsp_data <= 32'h275A7640;
        16'h1EC3C : rd_rsp_data <= 32'h05FC11C5;
        16'h1EC40 : rd_rsp_data <= 32'h28000600;
        16'h1EC44 : rd_rsp_data <= 32'h00004000;
        16'h1EC48 : rd_rsp_data <= 32'h00013880;
        16'h1EC4C : rd_rsp_data <= 32'h000004B3;
        16'h1EC50 : rd_rsp_data <= 32'h00000012;
        16'h1EC54 : rd_rsp_data <= 32'h00000001;
        16'h1EC58 : rd_rsp_data <= 32'h00001C00;
        16'h1EC6C : rd_rsp_data <= 32'h00000101;
        16'h1EC70 : rd_rsp_data <= 32'h00000101;
        16'h1EC74 : rd_rsp_data <= 32'h00422C80;
        16'h1EC78 : rd_rsp_data <= 32'h00000004;
        16'h1EC80 : rd_rsp_data <= 32'h23444688;
        16'h1EC88 : rd_rsp_data <= 32'h0AC4DC14;
        16'h1EC94 : rd_rsp_data <= 32'h11311022;
        16'h1EC98 : rd_rsp_data <= 32'h23444688;
        16'h1EC9C : rd_rsp_data <= 32'h00000008;
        16'h1ECB0 : rd_rsp_data <= 32'h0DC91596;
        16'h1ECB8 : rd_rsp_data <= 32'h23444688;
        16'h1ECBC : rd_rsp_data <= 32'h00000012;
        16'h1ECC0 : rd_rsp_data <= 32'h000002C2;
        16'h1ECC4 : rd_rsp_data <= 32'h02000140;
        16'h1ECC8 : rd_rsp_data <= 32'h0C078000;
        16'h1ECFC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1EDCC : rd_rsp_data <= 32'h3F000000;
        16'h1EDD0 : rd_rsp_data <= 32'hE0400000;
        16'h1EDD4 : rd_rsp_data <= 32'h26000400;
        16'h1EDE0 : rd_rsp_data <= 32'h00002003;
        16'h1EDE4 : rd_rsp_data <= 32'h0000000F;
        16'h1EDFC : rd_rsp_data <= 32'h08041000;
        16'h1EE00 : rd_rsp_data <= 32'h80400000;
        16'h1EE04 : rd_rsp_data <= 32'h8040010E;
        16'h1EE08 : rd_rsp_data <= 32'h80400201;
        16'h1EE0C : rd_rsp_data <= 32'h80400302;
        16'h1EE10 : rd_rsp_data <= 32'h80400405;
        16'h1EE14 : rd_rsp_data <= 32'h80400503;
        16'h1EE18 : rd_rsp_data <= 32'h80400604;
        16'h1EE1C : rd_rsp_data <= 32'h80400707;
        16'h1EE20 : rd_rsp_data <= 32'h8480080B;
        16'h1EE24 : rd_rsp_data <= 32'h8480090C;
        16'h1EE28 : rd_rsp_data <= 32'h80400A06;
        16'h1EE2C : rd_rsp_data <= 32'h80400B08;
        16'h1EE30 : rd_rsp_data <= 32'h80000C00;
        16'h1EE34 : rd_rsp_data <= 32'h80000D02;
        16'h1EE38 : rd_rsp_data <= 32'h80000E04;
        16'h1EE3C : rd_rsp_data <= 32'h80000F05;
        16'h1EE40 : rd_rsp_data <= 32'h80001006;
        16'h1EE44 : rd_rsp_data <= 32'h80001108;
        16'h1EE48 : rd_rsp_data <= 32'h8000120D;
        16'h1EE4C : rd_rsp_data <= 32'h8000130E;
        16'h1EE50 : rd_rsp_data <= 32'h80001481;
        16'h1EE54 : rd_rsp_data <= 32'h80001582;
        16'h1EE58 : rd_rsp_data <= 32'h80001683;
        16'h1EE5C : rd_rsp_data <= 32'h80001784;
        16'h1EE60 : rd_rsp_data <= 32'h80001489;
        16'h1EE64 : rd_rsp_data <= 32'h8000158A;
        16'h1EE68 : rd_rsp_data <= 32'h8000168B;
        16'h1EE6C : rd_rsp_data <= 32'h8000178C;
        16'h1EE70 : rd_rsp_data <= 32'h80001491;
        16'h1EE74 : rd_rsp_data <= 32'h80001592;
        16'h1EE78 : rd_rsp_data <= 32'h80001693;
        16'h1EE7C : rd_rsp_data <= 32'h80001794;
        16'h1EE80 : rd_rsp_data <= 32'h80001499;
        16'h1EE84 : rd_rsp_data <= 32'h8000159A;
        16'h1EE88 : rd_rsp_data <= 32'h8000169B;
        16'h1EE8C : rd_rsp_data <= 32'h8000179C;
        16'h1EE90 : rd_rsp_data <= 32'h800014A1;
        16'h1EE94 : rd_rsp_data <= 32'h800015A2;
        16'h1EE98 : rd_rsp_data <= 32'h800016A3;
        16'h1EE9C : rd_rsp_data <= 32'h800017A4;
        16'h1EEA0 : rd_rsp_data <= 32'h800014A9;
        16'h1EEA4 : rd_rsp_data <= 32'h800015AA;
        16'h1EEA8 : rd_rsp_data <= 32'h800016AB;
        16'h1EEAC : rd_rsp_data <= 32'h800017AC;
        16'h1EEB0 : rd_rsp_data <= 32'h800014B1;
        16'h1EEB4 : rd_rsp_data <= 32'h800015B2;
        16'h1EEB8 : rd_rsp_data <= 32'h800016B3;
        16'h1EEBC : rd_rsp_data <= 32'h800017B4;
        16'h1EEC0 : rd_rsp_data <= 32'h800014B9;
        16'h1EEC4 : rd_rsp_data <= 32'h800015BA;
        16'h1EEC8 : rd_rsp_data <= 32'h800016BB;
        16'h1EECC : rd_rsp_data <= 32'h800017BC;
        16'h1EED0 : rd_rsp_data <= 32'h800014C1;
        16'h1EED4 : rd_rsp_data <= 32'h800015C2;
        16'h1EED8 : rd_rsp_data <= 32'h800016C3;
        16'h1EEDC : rd_rsp_data <= 32'h800017C4;
        16'h1EEE0 : rd_rsp_data <= 32'h800014C9;
        16'h1EEE4 : rd_rsp_data <= 32'h800015CA;
        16'h1EEE8 : rd_rsp_data <= 32'h800016CB;
        16'h1EEEC : rd_rsp_data <= 32'h800017CC;
        16'h1EEF0 : rd_rsp_data <= 32'h800014D1;
        16'h1EEF4 : rd_rsp_data <= 32'h800015D2;
        16'h1EEF8 : rd_rsp_data <= 32'h800016D3;
        16'h1EEFC : rd_rsp_data <= 32'h800017D4;
        16'h1EF00 : rd_rsp_data <= 32'h800014D9;
        16'h1EF04 : rd_rsp_data <= 32'h800015DA;
        16'h1EF08 : rd_rsp_data <= 32'h800016DB;
        16'h1EF0C : rd_rsp_data <= 32'h800017DC;
        16'h1EF10 : rd_rsp_data <= 32'h800014E1;
        16'h1EF14 : rd_rsp_data <= 32'h800015E2;
        16'h1EF18 : rd_rsp_data <= 32'h800016E3;
        16'h1EF1C : rd_rsp_data <= 32'h800017E4;
        16'h1EF20 : rd_rsp_data <= 32'h800014E9;
        16'h1EF24 : rd_rsp_data <= 32'h800015EA;
        16'h1EF28 : rd_rsp_data <= 32'h800016EB;
        16'h1EF2C : rd_rsp_data <= 32'h800017EC;
        16'h1EF30 : rd_rsp_data <= 32'h800014F1;
        16'h1EF34 : rd_rsp_data <= 32'h800015F2;
        16'h1EF38 : rd_rsp_data <= 32'h800016F3;
        16'h1EF3C : rd_rsp_data <= 32'h800017F4;
        16'h1EF40 : rd_rsp_data <= 32'h800014F9;
        16'h1EF44 : rd_rsp_data <= 32'h800015FA;
        16'h1EF48 : rd_rsp_data <= 32'h800016FB;
        16'h1EF4C : rd_rsp_data <= 32'h830017FC;
        16'h1EF50 : rd_rsp_data <= 32'h80001822;
        16'h1EF54 : rd_rsp_data <= 32'h80001923;
        16'h1EF58 : rd_rsp_data <= 32'h80001A24;
        16'h1EF5C : rd_rsp_data <= 32'h80001B25;
        16'h1EF60 : rd_rsp_data <= 32'h80001C26;
        16'h1EF64 : rd_rsp_data <= 32'h80001D27;
        16'h1EF68 : rd_rsp_data <= 32'h80001E28;
        16'h1EF6C : rd_rsp_data <= 32'h80001F2D;
        16'h1EF70 : rd_rsp_data <= 32'hC800200A;
        16'h1EF74 : rd_rsp_data <= 32'hC8002203;
        16'h1EF78 : rd_rsp_data <= 32'h8040240F;
        16'h1F000 : rd_rsp_data <= 32'h27422027;
        16'h1F004 : rd_rsp_data <= 32'h01393075;
        16'h1F008 : rd_rsp_data <= 32'h49041828;
        16'h1F00C : rd_rsp_data <= 32'h0E0E088C;
        16'h1F010 : rd_rsp_data <= 32'h16141212;
        16'h1F014 : rd_rsp_data <= 32'h18306C48;
        16'h1F018 : rd_rsp_data <= 32'h0E0E081A;
        16'h1F01C : rd_rsp_data <= 32'h003FF020;
        16'h1F020 : rd_rsp_data <= 32'h19191944;
        16'h1F024 : rd_rsp_data <= 32'h19191919;
        16'h1F028 : rd_rsp_data <= 32'h80000020;
        16'h1F02C : rd_rsp_data <= 32'h4E000200;
        16'h1F034 : rd_rsp_data <= 32'h06010198;
        16'h1F038 : rd_rsp_data <= 32'h00000C00;
        16'h1F040 : rd_rsp_data <= 32'h00020208;
        16'h1F044 : rd_rsp_data <= 32'h00000200;
        16'h1F050 : rd_rsp_data <= 32'h060E8912;
        16'h1F054 : rd_rsp_data <= 32'h12068076;
        16'h1F068 : rd_rsp_data <= 32'h103B2838;
        16'h1F06C : rd_rsp_data <= 32'h16404030;
        16'h1F070 : rd_rsp_data <= 32'h26280000;
        16'h1F074 : rd_rsp_data <= 32'h00000080;
        16'h1F078 : rd_rsp_data <= 32'h00300004;
        16'h1F088 : rd_rsp_data <= 32'h8FC00029;
        16'h1F08C : rd_rsp_data <= 32'h0C008484;
        16'h1F090 : rd_rsp_data <= 32'h0C180810;
        16'h1F094 : rd_rsp_data <= 32'h08100408;
        16'h1F098 : rd_rsp_data <= 32'h040C0206;
        16'h1F0A0 : rd_rsp_data <= 32'hD4CA450A;
        16'h1F0A8 : rd_rsp_data <= 32'h02540040;
        16'h1F0AC : rd_rsp_data <= 32'h0281284B;
        16'h1F0B0 : rd_rsp_data <= 32'h0000000F;
        16'h1F0B8 : rd_rsp_data <= 32'h08104426;
        16'h1F0C0 : rd_rsp_data <= 32'h00200086;
        16'h1F0C4 : rd_rsp_data <= 32'h800308E2;
        16'h1F0C8 : rd_rsp_data <= 32'h1C483616;
        16'h1F0D0 : rd_rsp_data <= 32'h0000000F;
        16'h1F0D4 : rd_rsp_data <= 32'h0E64E893;
        16'h1F100 : rd_rsp_data <= 32'h80202028;
        16'h1F110 : rd_rsp_data <= 32'h00000056;
        16'h1F114 : rd_rsp_data <= 32'h00020611;
        16'h1F118 : rd_rsp_data <= 32'hFFF080AE;
        16'h1F11C : rd_rsp_data <= 32'h0001B20A;
        16'h1F120 : rd_rsp_data <= 32'h000000E0;
        16'h1F124 : rd_rsp_data <= 32'h00004000;
        16'h1F128 : rd_rsp_data <= 32'h20000000;
        16'h1F12C : rd_rsp_data <= 32'h00000007;
        16'h1F200 : rd_rsp_data <= 32'h30200884;
        16'h1F204 : rd_rsp_data <= 32'h4F3F2F40;
        16'h1F208 : rd_rsp_data <= 32'h5E56B733;
        16'h1F20C : rd_rsp_data <= 32'h00129024;
        16'h1F210 : rd_rsp_data <= 32'h00040844;
        16'h1F214 : rd_rsp_data <= 32'h80C3C3E8;
        16'h1F218 : rd_rsp_data <= 32'h1B000036;
        16'h1F21C : rd_rsp_data <= 32'h3F001B1B;
        16'h1F220 : rd_rsp_data <= 32'h33333939;
        16'h1F224 : rd_rsp_data <= 32'h0000007F;
        16'h1F3E0 : rd_rsp_data <= 32'h013E9828;
        16'h1F3E4 : rd_rsp_data <= 32'h0000508D;
        16'h1F3F0 : rd_rsp_data <= 32'hCA02BCBE;
        16'h1F3F4 : rd_rsp_data <= 32'hD90F74E9;
        16'h1F400 : rd_rsp_data <= 32'h11002EC3;
        16'h1F404 : rd_rsp_data <= 32'h0000000F;
        16'h1F40C : rd_rsp_data <= 32'h00000137;
        16'h1F410 : rd_rsp_data <= 32'h00200D05;
        16'h1F418 : rd_rsp_data <= 32'h02020202;
        16'h1F424 : rd_rsp_data <= 32'h00000001;
        16'h1F428 : rd_rsp_data <= 32'h01010101;
        16'h1F42C : rd_rsp_data <= 32'h00101020;
        16'h1F430 : rd_rsp_data <= 32'h23444688;
        16'h1F434 : rd_rsp_data <= 32'h00000008;
        16'h1F438 : rd_rsp_data <= 32'h275A7640;
        16'h1F43C : rd_rsp_data <= 32'h05FC11C5;
        16'h1F440 : rd_rsp_data <= 32'h28000600;
        16'h1F444 : rd_rsp_data <= 32'h00004000;
        16'h1F448 : rd_rsp_data <= 32'h00013880;
        16'h1F44C : rd_rsp_data <= 32'h000004B3;
        16'h1F450 : rd_rsp_data <= 32'h00000012;
        16'h1F454 : rd_rsp_data <= 32'h00000001;
        16'h1F458 : rd_rsp_data <= 32'h00001C00;
        16'h1F46C : rd_rsp_data <= 32'h00000101;
        16'h1F470 : rd_rsp_data <= 32'h00000101;
        16'h1F474 : rd_rsp_data <= 32'h0084B9C0;
        16'h1F478 : rd_rsp_data <= 32'h00000003;
        16'h1F480 : rd_rsp_data <= 32'h23444688;
        16'h1F484 : rd_rsp_data <= 32'h00000009;
        16'h1F488 : rd_rsp_data <= 32'h0AC4DC14;
        16'h1F494 : rd_rsp_data <= 32'h11311022;
        16'h1F498 : rd_rsp_data <= 32'h23444688;
        16'h1F49C : rd_rsp_data <= 32'h00000008;
        16'h1F4B0 : rd_rsp_data <= 32'h0DC910CB;
        16'h1F4B8 : rd_rsp_data <= 32'h23444688;
        16'h1F4BC : rd_rsp_data <= 32'h0000001B;
        16'h1F4C0 : rd_rsp_data <= 32'h000002C2;
        16'h1F4C4 : rd_rsp_data <= 32'h02000140;
        16'h1F4C8 : rd_rsp_data <= 32'h0C078000;
        16'h1F4D8 : rd_rsp_data <= 32'h854653C3;
        16'h1F4DC : rd_rsp_data <= 32'h56ABF65C;
        16'h1F4FC : rd_rsp_data <= 32'hFFFFFFFF;
        16'h1F5CC : rd_rsp_data <= 32'h3F000000;
        16'h1F5D0 : rd_rsp_data <= 32'hE0400000;
        16'h1F5D4 : rd_rsp_data <= 32'h26000400;
        16'h1F5E0 : rd_rsp_data <= 32'h00002003;
        16'h1F5E4 : rd_rsp_data <= 32'h0000000F;
        16'h1F5FC : rd_rsp_data <= 32'h08041000;
        16'h1F600 : rd_rsp_data <= 32'h80400000;
        16'h1F604 : rd_rsp_data <= 32'h8040010E;
        16'h1F608 : rd_rsp_data <= 32'h80400201;
        16'h1F60C : rd_rsp_data <= 32'h80400302;
        16'h1F610 : rd_rsp_data <= 32'h80400405;
        16'h1F614 : rd_rsp_data <= 32'h80400503;
        16'h1F618 : rd_rsp_data <= 32'h80400604;
        16'h1F61C : rd_rsp_data <= 32'h80400707;
        16'h1F620 : rd_rsp_data <= 32'h8480080B;
        16'h1F624 : rd_rsp_data <= 32'h8480090C;
        16'h1F628 : rd_rsp_data <= 32'h80400A06;
        16'h1F62C : rd_rsp_data <= 32'h80400B08;
        16'h1F630 : rd_rsp_data <= 32'h80000C00;
        16'h1F634 : rd_rsp_data <= 32'h80000D02;
        16'h1F638 : rd_rsp_data <= 32'h80000E04;
        16'h1F63C : rd_rsp_data <= 32'h80000F05;
        16'h1F640 : rd_rsp_data <= 32'h80001006;
        16'h1F644 : rd_rsp_data <= 32'h80001108;
        16'h1F648 : rd_rsp_data <= 32'h8000120D;
        16'h1F64C : rd_rsp_data <= 32'h8000130E;
        16'h1F650 : rd_rsp_data <= 32'h80001481;
        16'h1F654 : rd_rsp_data <= 32'h80001582;
        16'h1F658 : rd_rsp_data <= 32'h80001683;
        16'h1F65C : rd_rsp_data <= 32'h80001784;
        16'h1F660 : rd_rsp_data <= 32'h80001489;
        16'h1F664 : rd_rsp_data <= 32'h8000158A;
        16'h1F668 : rd_rsp_data <= 32'h8000168B;
        16'h1F66C : rd_rsp_data <= 32'h8000178C;
        16'h1F670 : rd_rsp_data <= 32'h80001491;
        16'h1F674 : rd_rsp_data <= 32'h80001592;
        16'h1F678 : rd_rsp_data <= 32'h80001693;
        16'h1F67C : rd_rsp_data <= 32'h80001794;
        16'h1F680 : rd_rsp_data <= 32'h80001499;
        16'h1F684 : rd_rsp_data <= 32'h8000159A;
        16'h1F688 : rd_rsp_data <= 32'h8000169B;
        16'h1F68C : rd_rsp_data <= 32'h8000179C;
        16'h1F690 : rd_rsp_data <= 32'h800014A1;
        16'h1F694 : rd_rsp_data <= 32'h800015A2;
        16'h1F698 : rd_rsp_data <= 32'h800016A3;
        16'h1F69C : rd_rsp_data <= 32'h800017A4;
        16'h1F6A0 : rd_rsp_data <= 32'h800014A9;
        16'h1F6A4 : rd_rsp_data <= 32'h800015AA;
        16'h1F6A8 : rd_rsp_data <= 32'h800016AB;
        16'h1F6AC : rd_rsp_data <= 32'h800017AC;
        16'h1F6B0 : rd_rsp_data <= 32'h800014B1;
        16'h1F6B4 : rd_rsp_data <= 32'h800015B2;
        16'h1F6B8 : rd_rsp_data <= 32'h800016B3;
        16'h1F6BC : rd_rsp_data <= 32'h800017B4;
        16'h1F6C0 : rd_rsp_data <= 32'h800014B9;
        16'h1F6C4 : rd_rsp_data <= 32'h800015BA;
        16'h1F6C8 : rd_rsp_data <= 32'h800016BB;
        16'h1F6CC : rd_rsp_data <= 32'h800017BC;
        16'h1F6D0 : rd_rsp_data <= 32'h800014C1;
        16'h1F6D4 : rd_rsp_data <= 32'h800015C2;
        16'h1F6D8 : rd_rsp_data <= 32'h800016C3;
        16'h1F6DC : rd_rsp_data <= 32'h800017C4;
        16'h1F6E0 : rd_rsp_data <= 32'h800014C9;
        16'h1F6E4 : rd_rsp_data <= 32'h800015CA;
        16'h1F6E8 : rd_rsp_data <= 32'h800016CB;
        16'h1F6EC : rd_rsp_data <= 32'h800017CC;
        16'h1F6F0 : rd_rsp_data <= 32'h800014D1;
        16'h1F6F4 : rd_rsp_data <= 32'h800015D2;
        16'h1F6F8 : rd_rsp_data <= 32'h800016D3;
        16'h1F6FC : rd_rsp_data <= 32'h800017D4;
        16'h1F700 : rd_rsp_data <= 32'h800014D9;
        16'h1F704 : rd_rsp_data <= 32'h800015DA;
        16'h1F708 : rd_rsp_data <= 32'h800016DB;
        16'h1F70C : rd_rsp_data <= 32'h800017DC;
        16'h1F710 : rd_rsp_data <= 32'h800014E1;
        16'h1F714 : rd_rsp_data <= 32'h800015E2;
        16'h1F718 : rd_rsp_data <= 32'h800016E3;
        16'h1F71C : rd_rsp_data <= 32'h800017E4;
        16'h1F720 : rd_rsp_data <= 32'h800014E9;
        16'h1F724 : rd_rsp_data <= 32'h800015EA;
        16'h1F728 : rd_rsp_data <= 32'h800016EB;
        16'h1F72C : rd_rsp_data <= 32'h800017EC;
        16'h1F730 : rd_rsp_data <= 32'h800014F1;
        16'h1F734 : rd_rsp_data <= 32'h800015F2;
        16'h1F738 : rd_rsp_data <= 32'h800016F3;
        16'h1F73C : rd_rsp_data <= 32'h800017F4;
        16'h1F740 : rd_rsp_data <= 32'h800014F9;
        16'h1F744 : rd_rsp_data <= 32'h800015FA;
        16'h1F748 : rd_rsp_data <= 32'h800016FB;
        16'h1F74C : rd_rsp_data <= 32'h830017FC;
        16'h1F750 : rd_rsp_data <= 32'h80001822;
        16'h1F754 : rd_rsp_data <= 32'h80001923;
        16'h1F758 : rd_rsp_data <= 32'h80001A24;
        16'h1F75C : rd_rsp_data <= 32'h80001B25;
        16'h1F760 : rd_rsp_data <= 32'h80001C26;
        16'h1F764 : rd_rsp_data <= 32'h80001D27;
        16'h1F768 : rd_rsp_data <= 32'h80001E28;
        16'h1F76C : rd_rsp_data <= 32'h80001F2D;
        16'h1F770 : rd_rsp_data <= 32'hC800200A;
        16'h1F774 : rd_rsp_data <= 32'hC8002203;
        16'h1F778 : rd_rsp_data <= 32'h8040240F;
        default: rd_rsp_data <= 32'h00000000;
    endcase
        end else if (dwr_valid) begin
            case (({dwr_addr[31:24], dwr_addr[23:16], dwr_addr[15:08], dwr_addr[07:00]}) & 32'hFFFFF)
            32'h599c : tj_max <= dwr_data;
            32'h597c : pp0_temp <= dwr_data;
            32'h5980 : pp1_temp <= dwr_data;
            32'h5978 : pkg_temp <= dwr_data;
            32'h5820 : thres <= dwr_data;
            32'h7200 : status <= dwr_data;
            endcase
        end else begin
            rd_rsp_data <= 32'h00000000;
        end
    end
            
endmodule



